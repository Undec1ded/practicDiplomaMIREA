`timescale 1ns / 1ps

//module for switching notes

module unravel#(
       
)(
    input clk,
    input button_action,
    
    output logic [3 : 0] note

);

reg [3 : 0] A1_note = 4'b0001;  //440
reg [3 : 0] Ah1_note = 4'b0010; //466 
reg [3 : 0] A2_note = 4'b0011;  //880
reg [3 : 0] Ah2_note = 4'b0100; //932
reg [3 : 0] C2_note = 4'b0101;  //523
reg [3 : 0] C3_note = 4'b0110;  //1046
reg [3 : 0] D2_note = 4'b0111;  //587
reg [3 : 0] Dh2_note = 4'b1000; //622
reg [3 : 0] D3_note = 4'b1001;  //1174
reg [3 : 0] F2_note = 4'b1010;  //698
reg [3 : 0] F3_note = 4'b1011;  //1396
reg [3 : 0] G1_note = 4'b1100;  //391
reg [3 : 0] G2_note = 4'b1101;  //783
reg [3 : 0] G3_note = 4'b1110;  //1567


reg [24 : 0] counter_sec = 0; 
reg [23 : 0] counter_time = 0;
reg time_driver = 0;
reg [3 : 0] state_note = 0;

//time_driver = 1 ms
always@ (posedge clk & counter_time != 100000) begin
    
    if (button_action == 1 & counter_time != 100000) begin
        time_driver = 0;
        counter_time = counter_time + 1;
    end
    else begin
        time_driver = 1;
        counter_time = 0;
end    
end

always@(posedge time_driver) begin
    if ((button_action) == 1) begin
        counter_sec = counter_sec + 1;
    end
    else begin 
        counter_sec = 0;
    end  
        case (counter_sec)
            0: note = Ah2_note;
            307: note = 0;
            341: note = C3_note;
            653: note = 0;
            688: note = Ah2_note;
            1000: note = 0;
            1035: note = Ah2_note;
            1191: note = 0;
            1209: note = G2_note;
            1365: note = 0;
            1556: note = C3_note;
            1868: note = 0;
            1903: note = Ah2_note;
            2215: note = 0;
            2250: note = A2_note;
            2562: note = 0;
            2597: note = G2_note;
            2909: note = 0;
            2944: note = G2_note;
            3100: note = 0;
            3118: note = F2_note;
            3274: note = 0;
            3639: note = F2_note;
            3795: note = 0;
            3813: note = Dh2_note;
            4125: note = 0;
            4160: note = F2_note;
            4316: note = 0;
            4334: note = D2_note;
            5115: note = 0;
            5723: note = D2_note;
            5879: note = 0;
            5897: note = D2_note;
            6209: note = 0;
            6244: note = D2_note;
            6400: note = 0;
            6418: note = D2_note;
            6730: note = 0;
            6765: note = C3_note;
            6921: note = 0;
            6939: note = C3_note;
            7251: note = 0;
            8501: note = Ah2_note;
            8657: note = 0;
            8675: note = A2_note;
            8987: note = 0;
            9022: note = A2_note;
            9178: note = 0;
            9196: note = A2_note;
            9508: note = 0;
            9543: note = Ah2_note;
            9855: note = 0;
            9890: note = Ah2_note;
            10202: note = 0;
            11278: note = Ah2_note;
            11434: note = 0;
            11452: note = C3_note;
            11764: note = 0;
            11799: note = Ah2_note;
            12111: note = 0;
            12146: note = A2_note;
            12302: note = 0;
            12320: note = G2_note;
            12476: note = 0;
            12667: note = C3_note;
            12979: note = 0;
            13014: note = Ah2_note;
            13326: note = 0;
            13361: note = A2_note;
            13673: note = 0;
            13708: note = G2_note;
            14020: note = 0;
            14055: note = G2_note;
            14211: note = 0;
            14229: note = F2_note;
            14541: note = 0;
            14749: note = F2_note;
            14905: note = 0;
            14923: note = Dh2_note;
            15235: note = 0;
            15270: note = F2_note;
            15426: note = 0;
            15444: note = D2_note;
            16068: note = 0;
            16833: note = D2_note;
            16989: note = 0;
            17007: note = D2_note;
            17319: note = 0;
            17354: note = D2_note;
            17510: note = 0;
            17528: note = D2_note;
            17840: note = 0;
            17875: note = C3_note;
            18031: note = 0;
            18049: note = C3_note;
            18361: note = 0;
            19611: note = Ah2_note;
            19767: note = 0;
            19785: note = A2_note;
            20097: note = 0;
            20132: note = A2_note;
            20288: note = 0;
            20306: note = A2_note;
            20618: note = 0;
            20653: note = Ah2_note;
            20965: note = 0;
            21000: note = Ah2_note;
            21156: note = 0;
            21174: note = D2_note;
            21251: note = 0;
            21261: note = D2_note;
            21338: note = 0;
            21435: note = D2_note;
            21512: note = 0;
            21609: note = D2_note;
            21686: note = 0;
            21696: note = D2_note;
            21773: note = 0;
            21870: note = D2_note;
            21947: note = 0;
            21957: note = D2_note;
            22034: note = 0;
            22131: note = D2_note;
            22208: note = 0;
            22305: note = D2_note;
            22382: note = 0;
            22392: note = D2_note;
            22469: note = 0;
            22566: note = D2_note;
            22643: note = 0;
            22653: note = G1_note;
            22730: note = 0;
            22740: note = G1_note;
            22817: note = 0;
            22827: note = A1_note;
            22904: note = 0;
            22914: note = G1_note;
            22991: note = 0;
            23001: note = G1_note;
            23078: note = 0;
            23088: note = Ah1_note;
            23165: note = 0;
            23175: note = A1_note;
            23252: note = 0;
            23262: note = D2_note;
            23339: note = 0;
            23349: note = G1_note;
            23426: note = 0;
            23436: note = G1_note;
            23513: note = 0;
            23523: note = A1_note;
            23600: note = 0;
            23610: note = G1_note;
            23687: note = 0;
            23697: note = G1_note;
            23774: note = 0;
            23784: note = A1_note;
            23861: note = 0;
            23871: note = G1_note;
            23948: note = 0;
            23958: note = D2_note;
            24035: note = 0;
            24045: note = D2_note;
            24122: note = 0;
            24219: note = D2_note;
            24296: note = 0;
            24393: note = D2_note;
            24470: note = 0;
            24480: note = D2_note;
            24557: note = 0;
            24654: note = D2_note;
            24731: note = 0;
            24741: note = D2_note;
            24818: note = 0;
            24915: note = D2_note;
            24992: note = 0;
            25089: note = D2_note;
            25166: note = 0;
            25176: note = D2_note;
            25253: note = 0;
            25350: note = D2_note;
            25427: note = 0;
            25437: note = Ah2_note;
            25514: note = 0;
            25611: note = D2_note;
            25688: note = 0;
            25698: note = G2_note;
            25854: note = 0;
            25872: note = Ah1_note;
            25949: note = 0;
            25959: note = Ah1_note;
            26036: note = 0;
            26046: note = C2_note;
            26123: note = 0;
            26133: note = Ah1_note;
            26210: note = 0;
            26220: note = G2_note;
            26297: note = 0;
            26307: note = Ah1_note;
            26384: note = 0;
            26394: note = Ah1_note;
            26471: note = 0;
            26481: note = F2_note;
            26558: note = 0;
            26568: note = Ah1_note;
            26724: note = 0;
            26742: note = Ah1_note;
            26819: note = 0;
            26829: note = Ah2_note;
            26906: note = 0;
            27003: note = D2_note;
            27080: note = 0;
            27090: note = G2_note;
            27246: note = 0;
            27264: note = Ah1_note;
            27341: note = 0;
            27351: note = Ah1_note;
            27428: note = 0;
            27438: note = C2_note;
            27515: note = 0;
            27525: note = Ah1_note;
            27602: note = 0;
            27612: note = G2_note;
            27689: note = 0;
            27699: note = Ah1_note;
            27776: note = 0;
            27786: note = Ah1_note;
            27863: note = 0;
            27873: note = G2_note;
            27950: note = 0;
            27960: note = Ah1_note;
            28116: note = 0;
            28134: note = Ah1_note;
            28211: note = 0;
            28221: note = Ah2_note;
            28298: note = 0;
            28395: note = D2_note;
            28472: note = 0;
            28482: note = G2_note;
            28638: note = 0;
            28656: note = Ah1_note;
            28733: note = 0;
            28743: note = Ah1_note;
            28820: note = 0;
            28830: note = C2_note;
            28907: note = 0;
            28917: note = Ah1_note;
            28994: note = 0;
            29004: note = G2_note;
            29081: note = 0;
            29091: note = Ah1_note;
            29168: note = 0;
            29178: note = Ah1_note;
            29255: note = 0;
            29265: note = G2_note;
            29342: note = 0;
            29352: note = Ah1_note;
            29508: note = 0;
            29526: note = Ah1_note;
            29603: note = 0;
            29613: note = Ah2_note;
            29690: note = 0;
            29787: note = D2_note;
            29864: note = 0;
            29874: note = G2_note;
            30030: note = 0;
            30048: note = Ah1_note;
            30125: note = 0;
            30135: note = Ah1_note;
            30212: note = 0;
            30222: note = C2_note;
            30299: note = 0;
            30309: note = Ah1_note;
            30386: note = 0;
            30396: note = G2_note;
            30473: note = 0;
            30483: note = Ah1_note;
            30560: note = 0;
            30570: note = Ah1_note;
            30647: note = 0;
            30657: note = G2_note;
            30734: note = 0;
            30744: note = Ah1_note;
            30900: note = 0;
            30918: note = F2_note;
            30995: note = 0;
            31005: note = G2_note;
            31082: note = 0;
            31179: note = Dh2_note;
            31256: note = 0;
            31439: note = A2_note;
            31516: note = 0;
            31613: note = F2_note;
            31690: note = 0;
            31700: note = G2_note;
            31777: note = 0;
            31874: note = Dh2_note;
            31951: note = 0;
            32134: note = A2_note;
            32290: note = 0;
            32308: note = Ah2_note;
            32542: note = 0;
            32569: note = Ah2_note;
            32803: note = 0;
            32830: note = Ah2_note;
            32986: note = 0;
            33351: note = Ah2_note;
            33507: note = 0;
            33525: note = D3_note;
            33681: note = 0;
            33699: note = D3_note;
            33933: note = 0;
            33960: note = C3_note;
            34194: note = 0;
            34221: note = C3_note;
            34377: note = 0;
            34916: note = Ah2_note;
            35072: note = 0;
            35090: note = C3_note;
            35324: note = 0;
            35351: note = Ah2_note;
            35585: note = 0;
            35612: note = A2_note;
            35924: note = 0;
            35959: note = F2_note;
            36271: note = 0;
            36306: note = D2_note;
            36462: note = 0;
            37695: note = A2_note;
            37851: note = 0;
            37869: note = Ah2_note;
            38025: note = 0;
            38043: note = Ah2_note;
            38120: note = 0;
            38130: note = Ah2_note;
            38442: note = 0;
            38737: note = Ah2_note;
            38893: note = 0;
            39084: note = D3_note;
            39240: note = 0;
            39258: note = D3_note;
            39492: note = 0;
            39519: note = C3_note;
            39753: note = 0;
            39780: note = C3_note;
            40092: note = 0;
            40127: note = Ah2_note;
            40283: note = 0;
            40648: note = D3_note;
            40960: note = 0;
            40995: note = C3_note;
            41151: note = 0;
            41169: note = C3_note;
            41637: note = 0;
            41690: note = A2_note;
            41846: note = 0;
            41864: note = Ah2_note;
            42020: note = 0;
            43253: note = F3_note;
            43409: note = 0;
            43427: note = F3_note;
            43583: note = 0;
            43601: note = D3_note;
            43678: note = 0;
            43688: note = D3_note;
            43765: note = 0;
            43948: note = D3_note;
            44104: note = 0;
            44122: note = C3_note;
            44278: note = 0;
            44296: note = D3_note;
            44373: note = 0;
            44383: note = D3_note;
            44460: note = 0;
            44643: note = F3_note;
            44799: note = 0;
            44817: note = F3_note;
            44973: note = 0;
            44991: note = D3_note;
            45068: note = 0;
            45078: note = D3_note;
            45155: note = 0;
            45338: note = D3_note;
            45494: note = 0;
            45512: note = C3_note;
            45668: note = 0;
            45686: note = D3_note;
            45763: note = 0;
            45773: note = D3_note;
            45850: note = 0;
            46033: note = F3_note;
            46189: note = 0;
            46207: note = F3_note;
            46363: note = 0;
            46381: note = D3_note;
            46458: note = 0;
            46468: note = D3_note;
            46545: note = 0;
            46728: note = D3_note;
            46884: note = 0;
            46902: note = C3_note;
            47136: note = 0;
            47163: note = C3_note;
            47397: note = 0;
            47424: note = C3_note;
            47580: note = 0;
            47598: note = D3_note;
            48066: note = 0;
            48119: note = D3_note;
            48275: note = 0;
            48293: note = D3_note;
            48527: note = 0;
            48554: note = C3_note;
            48788: note = 0;
            48815: note = C3_note;
            48971: note = 0;
            48989: note = D3_note;
            49223: note = 0;
            49250: note = C3_note;
            49484: note = 0;
            49511: note = C3_note;
            49667: note = 0;
            49685: note = C3_note;
            49919: note = 0;
            49946: note = Ah2_note;
            50180: note = 0;
            50207: note = Ah2_note;
            50363: note = 0;
            50381: note = A2_note;
            50615: note = 0;
            50642: note = Ah2_note;
            50876: note = 0;
            50903: note = A2_note;
            51215: note = 0;
            51250: note = F2_note;
            51562: note = 0;
            51597: note = F2_note;
            51753: note = 0;
            51771: note = D3_note;
            52005: note = 0;
            52032: note = C3_note;
            52266: note = 0;
            52293: note = C3_note;
            52449: note = 0;
            52467: note = C3_note;
            52701: note = 0;
            52728: note = Ah2_note;
            52962: note = 0;
            52989: note = Ah2_note;
            53145: note = 0;
            53163: note = A2_note;
            53397: note = 0;
            53424: note = Ah2_note;
            53658: note = 0;
            53685: note = F3_note;
            53997: note = 0;
            54032: note = A2_note;
            54344: note = 0;
            54379: note = A2_note;
            54535: note = 0;
            54553: note = G3_note;
            54787: note = 0;
            54814: note = F3_note;
            55048: note = 0;
            55075: note = F3_note;
            55231: note = 0;
            55249: note = F3_note;
            55483: note = 0;
            55510: note = D3_note;
            55744: note = 0;
            55771: note = Ah2_note;
            55927: note = 0;
            55945: note = Ah2_note;
            56179: note = 0;
            56206: note = A2_note;
            56440: note = 0;
            56467: note = G2_note;
            56779: note = 0;
            56814: note = A2_note;
            57126: note = 0;
            57161: note = Ah2_note;
            57785: note = 0;
            58550: note = Ah2_note;
            58706: note = 0;
            58724: note = A2_note;
            58958: note = 0;
            58985: note = Ah2_note;
            59219: note = 0;
            59246: note = A2_note;
            59558: note = 0;
            59593: note = F2_note;
            59905: note = 0;
            60113: note = D3_note;
            60347: note = 0;
            60374: note = C3_note;
            60608: note = 0;
            60635: note = C3_note;
            60791: note = 0;
            60809: note = C3_note;
            61043: note = 0;
            61070: note = Ah2_note;
            61304: note = 0;
            61331: note = Ah2_note;
            61487: note = 0;
            61505: note = A2_note;
            61739: note = 0;
            61766: note = Ah2_note;
            62000: note = 0;
            62027: note = A2_note;
            62339: note = 0;
            62374: note = F2_note;
            62686: note = 0;
            62721: note = F2_note;
            62877: note = 0;
            62895: note = D3_note;
            63129: note = 0;
            63156: note = C3_note;
            63390: note = 0;
            63417: note = C3_note;
            63573: note = 0;
            63591: note = C3_note;
            63825: note = 0;
            63852: note = Ah2_note;
            64086: note = 0;
            64113: note = Ah2_note;
            64269: note = 0;
            64287: note = A2_note;
            64521: note = 0;
            64548: note = Ah2_note;
            64782: note = 0;
            64809: note = F3_note;
            65121: note = 0;
            65156: note = A2_note;
            65468: note = 0;
            65503: note = A2_note;
            65659: note = 0;
            65677: note = G3_note;
            65911: note = 0;
            65938: note = F3_note;
            66172: note = 0;
            66199: note = F3_note;
            66355: note = 0;
            66373: note = F3_note;
            66607: note = 0;
            66634: note = D3_note;
            66868: note = 0;
            66895: note = Ah2_note;
            67051: note = 0;
            67069: note = Ah2_note;
            67303: note = 0;
            67330: note = A2_note;
            67564: note = 0;
            67591: note = G2_note;
            67903: note = 0;
            67938: note = A2_note;
            68250: note = 0;
            68285: note = Ah2_note;
            69691: note = 0;

        endcase  
end

endmodule