`timescale 1ns / 1ps

//module for switching notes

module unravel#(
       
)(
    input clk,
    input button_action,
    input [3 : 0] sw,
    
    output logic [5 : 0] note

);




reg [5 : 0] A1_note =  6'b000001;  //440
reg [5 : 0] Ah1_note = 6'b000010; //466 
reg [5 : 0] A2_note =  6'b000011;  //880
reg [5 : 0] Ah2_note = 6'b000100; //932
reg [5 : 0] C2_note = 6'b000101;  //523
reg [5 : 0] C3_note = 6'b000110;  //1046
reg [5 : 0] D2_note = 6'b000111;  //587
reg [5 : 0] F2_note = 6'b001010;  //698
reg [5 : 0] F3_note = 6'b001011;  //1396
reg [5 : 0] G1_note = 6'b001100;  //391
reg [5 : 0] G2_note = 6'b001101;  //783
reg [5 : 0] G3_note = 6'b001110;  //1567

reg [5 : 0] C1_note  = 6'b001111; //261
reg [5 : 0] Ch1_note = 6'b010000; //277
reg [5 : 0] Ch2_note = 6'b010001; //554
reg [5 : 0] Ch3_note = 6'b010010; //1108
reg [5 : 0] C4_note  = 6'b010011; //2093
reg [5 : 0] Ch4_note = 6'b010100; //2217
reg [5 : 0] D1_note  = 6'b010101; //293
reg [5 : 0] Dh1_note = 6'b010111; //311
reg [5 : 0] Dh2_note = 6'b011000; //622
reg [5 : 0] D3_note  = 6'b011001; //1174
reg [5 : 0] Dh3_note = 6'b011010; //1244
reg [5 : 0] D4_note  = 6'b011011; //2349
reg [5 : 0] Dh4_note = 6'b011100; //2489
reg [5 : 0] E1_note  = 6'b011101; //329
reg [5 : 0] E2_note  = 6'b011110; //659
reg [5 : 0] E3_note  = 6'b011111; //1318
reg [5 : 0] E4_note  = 6'b100000; //2637
reg [5 : 0] F1_note  = 6'b100001; //349
reg [5 : 0] Fh1_note = 6'b100010; //369
reg [5 : 0] Fh2_note = 6'b100011; //739
reg [5 : 0] Fh3_note = 6'b100101; //1480
reg [5 : 0] F4_note  = 6'b100110; //2793
reg [5 : 0] Fh4_note = 6'b100111; //2960
reg [5 : 0] Gh1_note = 6'b100111; //415
reg [5 : 0] Gh2_note = 6'b101000; //830
reg [5 : 0] Gh3_note = 6'b101001; //1661
reg [5 : 0] G4_note  = 6'b101010; //3136
reg [5 : 0] Gh4_note = 6'b101011; //3332
reg [5 : 0] A3_note  = 6'b101100; //1720
reg [5 : 0] Ah3_note = 6'b101101; //1864
reg [5 : 0] A4_note  = 6'b101110; //3440
reg [5 : 0] Ah4_note = 6'b101111; //3729
reg [5 : 0] B1_note  = 6'b110000; //493
reg [5 : 0] B2_note  = 6'b110001; //987
reg [5 : 0] B3_note  = 6'b110010; //1975
reg [5 : 0] B4_note  = 6'b110011; //3951
reg [5 : 0] C_note   = 6'b110100; //130
reg [5 : 0] Ch_note  = 6'b110101; //138
reg [5 : 0] D_note   = 6'b110110; //147
reg [5 : 0] Dh_note  = 6'b110111; //155
reg [5 : 0] E_note   = 6'b111000; //164
reg [5 : 0] F_note   = 6'b111001; //174
reg [5 : 0] Fh_note  = 6'b111010; //185
reg [5 : 0] G_note   = 6'b111011; //196
reg [5 : 0] Gh_note  = 6'b111100; //207
reg [5 : 0] A_note   = 6'b111101; //220
reg [5 : 0] Ah_note  = 6'b111110; //233
reg [5 : 0] B_note   = 6'b111111; //246

reg [24 : 0] counter_sec = 0; 
reg [23 : 0] counter_time = 0;
reg time_driver = 0;
reg [3 : 0] sw_state = 0;
//time_driver = 1 ms
always@ (posedge clk) begin
    sw_state = {sw[3], sw[2], sw[1], sw[0]};
    if (button_action == 1 & counter_time != 100000) begin
        time_driver = 0;
        counter_time = counter_time + 1;
    end
    else begin
        time_driver = 1;
        counter_time = 0;
end    
end

always@(posedge time_driver) begin
    if ((button_action) == 1) begin
        counter_sec = counter_sec + 1;
    end
    else begin 
        counter_sec = 0;
    end  
    //unravel
    if (sw_state == 4'b0001) begin
        case (counter_sec)
            2: note = Ah2_note;
            307: note = 0;
            341: note = C3_note;
            653: note = 0;
            688: note = Ah2_note;
            1000: note = 0;
            1035: note = Ah2_note;
            1191: note = 0;
            1209: note = G2_note;
            1365: note = 0;
            1556: note = C3_note;
            1868: note = 0;
            1903: note = Ah2_note;
            2215: note = 0;
            2250: note = A2_note;
            2562: note = 0;
            2597: note = G2_note;
            2909: note = 0;
            2944: note = G2_note;
            3100: note = 0;
            3118: note = F2_note;
            3274: note = 0;
            3639: note = F2_note;
            3795: note = 0;
            3813: note = Dh2_note;
            4125: note = 0;
            4160: note = F2_note;
            4316: note = 0;
            4334: note = D2_note;
            5115: note = 0;
            5723: note = D2_note;
            5879: note = 0;
            5897: note = D2_note;
            6209: note = 0;
            6244: note = D2_note;
            6400: note = 0;
            6418: note = D2_note;
            6730: note = 0;
            6765: note = C3_note;
            6921: note = 0;
            6939: note = C3_note;
            7251: note = 0;
            8501: note = Ah2_note;
            8657: note = 0;
            8675: note = A2_note;
            8987: note = 0;
            9022: note = A2_note;
            9178: note = 0;
            9196: note = A2_note;
            9508: note = 0;
            9543: note = Ah2_note;
            9855: note = 0;
            9890: note = Ah2_note;
            10202: note = 0;
            11278: note = Ah2_note;
            11434: note = 0;
            11452: note = C3_note;
            11764: note = 0;
            11799: note = Ah2_note;
            12111: note = 0;
            12146: note = A2_note;
            12302: note = 0;
            12320: note = G2_note;
            12476: note = 0;
            12667: note = C3_note;
            12979: note = 0;
            13014: note = Ah2_note;
            13326: note = 0;
            13361: note = A2_note;
            13673: note = 0;
            13708: note = G2_note;
            14020: note = 0;
            14055: note = G2_note;
            14211: note = 0;
            14229: note = F2_note;
            14541: note = 0;
            14749: note = F2_note;
            14905: note = 0;
            14923: note = Dh2_note;
            15235: note = 0;
            15270: note = F2_note;
            15426: note = 0;
            15444: note = D2_note;
            16068: note = 0;
            16833: note = D2_note;
            16989: note = 0;
            17007: note = D2_note;
            17319: note = 0;
            17354: note = D2_note;
            17510: note = 0;
            17528: note = D2_note;
            17840: note = 0;
            17875: note = C3_note;
            18031: note = 0;
            18049: note = C3_note;
            18361: note = 0;
            19611: note = Ah2_note;
            19767: note = 0;
            19785: note = A2_note;
            20097: note = 0;
            20132: note = A2_note;
            20288: note = 0;
            20306: note = A2_note;
            20618: note = 0;
            20653: note = Ah2_note;
            20965: note = 0;
            21000: note = Ah2_note;
            21156: note = 0;
            21174: note = D2_note;
            21251: note = 0;
            21261: note = D2_note;
            21338: note = 0;
            21435: note = D2_note;
            21512: note = 0;
            21609: note = D2_note;
            21686: note = 0;
            21696: note = D2_note;
            21773: note = 0;
            21870: note = D2_note;
            21947: note = 0;
            21957: note = D2_note;
            22034: note = 0;
            22131: note = D2_note;
            22208: note = 0;
            22305: note = D2_note;
            22382: note = 0;
            22392: note = D2_note;
            22469: note = 0;
            22566: note = D2_note;
            22643: note = 0;
            22653: note = G1_note;
            22730: note = 0;
            22740: note = G1_note;
            22817: note = 0;
            22827: note = A1_note;
            22904: note = 0;
            22914: note = G1_note;
            22991: note = 0;
            23001: note = G1_note;
            23078: note = 0;
            23088: note = Ah1_note;
            23165: note = 0;
            23175: note = A1_note;
            23252: note = 0;
            23262: note = D2_note;
            23339: note = 0;
            23349: note = G1_note;
            23426: note = 0;
            23436: note = G1_note;
            23513: note = 0;
            23523: note = A1_note;
            23600: note = 0;
            23610: note = G1_note;
            23687: note = 0;
            23697: note = G1_note;
            23774: note = 0;
            23784: note = A1_note;
            23861: note = 0;
            23871: note = G1_note;
            23948: note = 0;
            23958: note = D2_note;
            24035: note = 0;
            24045: note = D2_note;
            24122: note = 0;
            24219: note = D2_note;
            24296: note = 0;
            24393: note = D2_note;
            24470: note = 0;
            24480: note = D2_note;
            24557: note = 0;
            24654: note = D2_note;
            24731: note = 0;
            24741: note = D2_note;
            24818: note = 0;
            24915: note = D2_note;
            24992: note = 0;
            25089: note = D2_note;
            25166: note = 0;
            25176: note = D2_note;
            25253: note = 0;
            25350: note = D2_note;
            25427: note = 0;
            25437: note = Ah2_note;
            25514: note = 0;
            25611: note = D2_note;
            25688: note = 0;
            25698: note = G2_note;
            25854: note = 0;
            25872: note = Ah1_note;
            25949: note = 0;
            25959: note = Ah1_note;
            26036: note = 0;
            26046: note = C2_note;
            26123: note = 0;
            26133: note = Ah1_note;
            26210: note = 0;
            26220: note = G2_note;
            26297: note = 0;
            26307: note = Ah1_note;
            26384: note = 0;
            26394: note = Ah1_note;
            26471: note = 0;
            26481: note = F2_note;
            26558: note = 0;
            26568: note = Ah1_note;
            26724: note = 0;
            26742: note = Ah1_note;
            26819: note = 0;
            26829: note = Ah2_note;
            26906: note = 0;
            27003: note = D2_note;
            27080: note = 0;
            27090: note = G2_note;
            27246: note = 0;
            27264: note = Ah1_note;
            27341: note = 0;
            27351: note = Ah1_note;
            27428: note = 0;
            27438: note = C2_note;
            27515: note = 0;
            27525: note = Ah1_note;
            27602: note = 0;
            27612: note = G2_note;
            27689: note = 0;
            27699: note = Ah1_note;
            27776: note = 0;
            27786: note = Ah1_note;
            27863: note = 0;
            27873: note = G2_note;
            27950: note = 0;
            27960: note = Ah1_note;
            28116: note = 0;
            28134: note = Ah1_note;
            28211: note = 0;
            28221: note = Ah2_note;
            28298: note = 0;
            28395: note = D2_note;
            28472: note = 0;
            28482: note = G2_note;
            28638: note = 0;
            28656: note = Ah1_note;
            28733: note = 0;
            28743: note = Ah1_note;
            28820: note = 0;
            28830: note = C2_note;
            28907: note = 0;
            28917: note = Ah1_note;
            28994: note = 0;
            29004: note = G2_note;
            29081: note = 0;
            29091: note = Ah1_note;
            29168: note = 0;
            29178: note = Ah1_note;
            29255: note = 0;
            29265: note = G2_note;
            29342: note = 0;
            29352: note = Ah1_note;
            29508: note = 0;
            29526: note = Ah1_note;
            29603: note = 0;
            29613: note = Ah2_note;
            29690: note = 0;
            29787: note = D2_note;
            29864: note = 0;
            29874: note = G2_note;
            30030: note = 0;
            30048: note = Ah1_note;
            30125: note = 0;
            30135: note = Ah1_note;
            30212: note = 0;
            30222: note = C2_note;
            30299: note = 0;
            30309: note = Ah1_note;
            30386: note = 0;
            30396: note = G2_note;
            30473: note = 0;
            30483: note = Ah1_note;
            30560: note = 0;
            30570: note = Ah1_note;
            30647: note = 0;
            30657: note = G2_note;
            30734: note = 0;
            30744: note = Ah1_note;
            30900: note = 0;
            30918: note = F2_note;
            30995: note = 0;
            31005: note = G2_note;
            31082: note = 0;
            31179: note = Dh2_note;
            31256: note = 0;
            31439: note = A2_note;
            31516: note = 0;
            31613: note = F2_note;
            31690: note = 0;
            31700: note = G2_note;
            31777: note = 0;
            31874: note = Dh2_note;
            31951: note = 0;
            32134: note = A2_note;
            32290: note = 0;
            32308: note = Ah2_note;
            32542: note = 0;
            32569: note = Ah2_note;
            32803: note = 0;
            32830: note = Ah2_note;
            32986: note = 0;
            33351: note = Ah2_note;
            33507: note = 0;
            33525: note = D3_note;
            33681: note = 0;
            33699: note = D3_note;
            33933: note = 0;
            33960: note = C3_note;
            34194: note = 0;
            34221: note = C3_note;
            34377: note = 0;
            34916: note = Ah2_note;
            35072: note = 0;
            35090: note = C3_note;
            35324: note = 0;
            35351: note = Ah2_note;
            35585: note = 0;
            35612: note = A2_note;
            35924: note = 0;
            35959: note = F2_note;
            36271: note = 0;
            36306: note = D2_note;
            36462: note = 0;
            37695: note = A2_note;
            37851: note = 0;
            37869: note = Ah2_note;
            38025: note = 0;
            38043: note = Ah2_note;
            38120: note = 0;
            38130: note = Ah2_note;
            38442: note = 0;
            38737: note = Ah2_note;
            38893: note = 0;
            39084: note = D3_note;
            39240: note = 0;
            39258: note = D3_note;
            39492: note = 0;
            39519: note = C3_note;
            39753: note = 0;
            39780: note = C3_note;
            40092: note = 0;
            40127: note = Ah2_note;
            40283: note = 0;
            40648: note = D3_note;
            40960: note = 0;
            40995: note = C3_note;
            41151: note = 0;
            41169: note = C3_note;
            41637: note = 0;
            41690: note = A2_note;
            41846: note = 0;
            41864: note = Ah2_note;
            42020: note = 0;
            43253: note = F3_note;
            43409: note = 0;
            43427: note = F3_note;
            43583: note = 0;
            43601: note = D3_note;
            43678: note = 0;
            43688: note = D3_note;
            43765: note = 0;
            43948: note = D3_note;
            44104: note = 0;
            44122: note = C3_note;
            44278: note = 0;
            44296: note = D3_note;
            44373: note = 0;
            44383: note = D3_note;
            44460: note = 0;
            44643: note = F3_note;
            44799: note = 0;
            44817: note = F3_note;
            44973: note = 0;
            44991: note = D3_note;
            45068: note = 0;
            45078: note = D3_note;
            45155: note = 0;
            45338: note = D3_note;
            45494: note = 0;
            45512: note = C3_note;
            45668: note = 0;
            45686: note = D3_note;
            45763: note = 0;
            45773: note = D3_note;
            45850: note = 0;
            46033: note = F3_note;
            46189: note = 0;
            46207: note = F3_note;
            46363: note = 0;
            46381: note = D3_note;
            46458: note = 0;
            46468: note = D3_note;
            46545: note = 0;
            46728: note = D3_note;
            46884: note = 0;
            46902: note = C3_note;
            47136: note = 0;
            47163: note = C3_note;
            47397: note = 0;
            47424: note = C3_note;
            47580: note = 0;
            47598: note = D3_note;
            48066: note = 0;
            48119: note = D3_note;
            48275: note = 0;
            48293: note = D3_note;
            48527: note = 0;
            48554: note = C3_note;
            48788: note = 0;
            48815: note = C3_note;
            48971: note = 0;
            48989: note = D3_note;
            49223: note = 0;
            49250: note = C3_note;
            49484: note = 0;
            49511: note = C3_note;
            49667: note = 0;
            49685: note = C3_note;
            49919: note = 0;
            49946: note = Ah2_note;
            50180: note = 0;
            50207: note = Ah2_note;
            50363: note = 0;
            50381: note = A2_note;
            50615: note = 0;
            50642: note = Ah2_note;
            50876: note = 0;
            50903: note = A2_note;
            51215: note = 0;
            51250: note = F2_note;
            51562: note = 0;
            51597: note = F2_note;
            51753: note = 0;
            51771: note = D3_note;
            52005: note = 0;
            52032: note = C3_note;
            52266: note = 0;
            52293: note = C3_note;
            52449: note = 0;
            52467: note = C3_note;
            52701: note = 0;
            52728: note = Ah2_note;
            52962: note = 0;
            52989: note = Ah2_note;
            53145: note = 0;
            53163: note = A2_note;
            53397: note = 0;
            53424: note = Ah2_note;
            53658: note = 0;
            53685: note = F3_note;
            53997: note = 0;
            54032: note = A2_note;
            54344: note = 0;
            54379: note = A2_note;
            54535: note = 0;
            54553: note = G3_note;
            54787: note = 0;
            54814: note = F3_note;
            55048: note = 0;
            55075: note = F3_note;
            55231: note = 0;
            55249: note = F3_note;
            55483: note = 0;
            55510: note = D3_note;
            55744: note = 0;
            55771: note = Ah2_note;
            55927: note = 0;
            55945: note = Ah2_note;
            56179: note = 0;
            56206: note = A2_note;
            56440: note = 0;
            56467: note = G2_note;
            56779: note = 0;
            56814: note = A2_note;
            57126: note = 0;
            57161: note = Ah2_note;
            57785: note = 0;
            58550: note = Ah2_note;
            58706: note = 0;
            58724: note = A2_note;
            58958: note = 0;
            58985: note = Ah2_note;
            59219: note = 0;
            59246: note = A2_note;
            59558: note = 0;
            59593: note = F2_note;
            59905: note = 0;
            60113: note = D3_note;
            60347: note = 0;
            60374: note = C3_note;
            60608: note = 0;
            60635: note = C3_note;
            60791: note = 0;
            60809: note = C3_note;
            61043: note = 0;
            61070: note = Ah2_note;
            61304: note = 0;
            61331: note = Ah2_note;
            61487: note = 0;
            61505: note = A2_note;
            61739: note = 0;
            61766: note = Ah2_note;
            62000: note = 0;
            62027: note = A2_note;
            62339: note = 0;
            62374: note = F2_note;
            62686: note = 0;
            62721: note = F2_note;
            62877: note = 0;
            62895: note = D3_note;
            63129: note = 0;
            63156: note = C3_note;
            63390: note = 0;
            63417: note = C3_note;
            63573: note = 0;
            63591: note = C3_note;
            63825: note = 0;
            63852: note = Ah2_note;
            64086: note = 0;
            64113: note = Ah2_note;
            64269: note = 0;
            64287: note = A2_note;
            64521: note = 0;
            64548: note = Ah2_note;
            64782: note = 0;
            64809: note = F3_note;
            65121: note = 0;
            65156: note = A2_note;
            65468: note = 0;
            65503: note = A2_note;
            65659: note = 0;
            65677: note = G3_note;
            65911: note = 0;
            65938: note = F3_note;
            66172: note = 0;
            66199: note = F3_note;
            66355: note = 0;
            66373: note = F3_note;
            66607: note = 0;
            66634: note = D3_note;
            66868: note = 0;
            66895: note = Ah2_note;
            67051: note = 0;
            67069: note = Ah2_note;
            67303: note = 0;
            67330: note = A2_note;
            67564: note = 0;
            67591: note = G2_note;
            67903: note = 0;
            67938: note = A2_note;
            68250: note = 0;
            68285: note = Ah2_note;
            69691: note = 0;

        endcase  
    end 
    //falling
    else if (sw_state == 4'b0010) begin
        case (counter_sec)
            2'b11: note = Ah1_note;
            9'b101010000: note = 0;
            9'b110001010: note = Ch2_note;
            10'b1011011010: note = 0;
            10'b1100010100: note = Ah1_note;
            10'b1110111100: note = 0;
            10'b1111011001: note = Ch2_note;
            11'b10010000001: note = 0;
            11'b10010011110: note = Ch2_note;
            11'b10111101110: note = 0;
            11'b11000101000: note = Ah1_note;
            11'b11101111000: note = 0;
            11'b11110110010: note = Ch2_note;
            12'b100100000010: note = 0;
            12'b100100111100: note = Ah1_note;
            12'b101010001100: note = 0;
            12'b101011000110: note = Ch2_note;
            12'b110000010110: note = 0;
            12'b110001010000: note = Ah1_note;
            12'b110110100000: note = 0;
            12'b110111011010: note = Ch2_note;
            12'b111100101010: note = 0;
            12'b111101100100: note = Ah1_note;
            13'b1000000001100: note = 0;
            13'b1000000101001: note = Ch2_note;
            13'b1000011010001: note = 0;
            13'b1000011101110: note = Ch2_note;
            13'b1001000111110: note = 0;
            13'b1001100111100: note = Ch2_note;
            13'b1001111100100: note = 0;
            13'b1010000000001: note = Ch2_note;
            13'b1010101010001: note = 0;
            13'b1010110001011: note = Ah1_note;
            13'b1011000110011: note = 0;
            13'b1011001010000: note = Ch2_note;
            13'b1011011111000: note = 0;
            13'b1011100010101: note = Ch2_note;
            13'b1100001100101: note = 0;
            13'b1100010011111: note = Ah1_note;
            13'b1100111101111: note = 0;
            13'b1101000101001: note = Ch2_note;
            13'b1101101111001: note = 0;
            13'b1101110110011: note = Ah1_note;
            13'b1110001011011: note = 0;
            13'b1110001111000: note = Ch2_note;
            13'b1110100100000: note = 0;
            13'b1110100111101: note = Ch2_note;
            13'b1110111100101: note = 0;
            13'b1111000000010: note = Dh2_note;
            13'b1111010101010: note = 0;
            13'b1111011000111: note = F2_note;
            14'b10000010111111: note = 0;
            14'b10000100010101: note = Gh2_note;
            14'b10000110111101: note = 0;
            14'b10000111011010: note = F2_note;
            14'b10001100101010: note = 0;
            14'b10001101100100: note = Dh2_note;
            14'b10010010110100: note = 0;
            14'b10010011101110: note = Ch2_note;
            14'b10011110001110: note = 0;
            14'b10100011000110: note = C3_note;
            14'b10100101101110: note = 0;
            14'b10100110001011: note = Ch3_note;
            14'b10101000110011: note = 0;
            14'b10101001010000: note = Dh3_note;
            14'b10101011111000: note = 0;
            14'b10101100010101: note = C3_note;
            14'b10110110110101: note = 0;
            14'b10111000101000: note = Ah1_note;
            14'b10111011010000: note = 0;
            14'b10111011101101: note = Ch2_note;
            14'b10111110010101: note = 0;
            14'b10111110110010: note = Ch2_note;
            14'b11000001011010: note = 0;
            14'b11000001110111: note = Ch1_note;
            14'b11000100011111: note = 0;
            14'b11000100111100: note = Ch1_note;
            14'b11001000011100: note = 0;
            14'b11001001000011: note = Ch1_note;
            14'b11001100100011: note = 0;
            14'b11001101001010: note = Ch1_note;
            14'b11010000101010: note = 0;
            14'b11010001010001: note = Ch1_note;
            14'b11010100110001: note = 0;
            14'b11010101011000: note = Ch1_note;
            14'b11011000111000: note = 0;
            14'b11011001011111: note = F1_note;
            14'b11011100111111: note = 0;
            14'b11011101100110: note = C1_note;
            14'b11100001000110: note = 0;
            14'b11100001101101: note = C1_note;
            14'b11100101001101: note = 0;
            14'b11100101110100: note = C1_note;
            14'b11101001010100: note = 0;
            14'b11101001111011: note = C1_note;
            14'b11101100100011: note = 0;
            14'b11101101000000: note = C1_note;
            14'b11101111101000: note = 0;
            14'b11110000000101: note = C1_note;
            14'b11110010101101: note = 0;
            14'b11110011001010: note = C1_note;
            14'b11110101110010: note = 0;
            14'b11110110001111: note = Ch1_note;
            14'b11111001101111: note = 0;
            14'b11111010010110: note = Ch1_note;
            14'b11111101110110: note = 0;
            14'b11111110011101: note = Ch1_note;
            15'b100000001111101: note = 0;
            15'b100000010100100: note = Ch1_note;
            15'b100000110000100: note = 0;
            15'b100000110101011: note = Ch1_note;
            15'b100001010001011: note = 0;
            15'b100001010110010: note = F1_note;
            15'b100001110010010: note = 0;
            15'b100001110111001: note = C1_note;
            15'b100010010011001: note = 0;
            15'b100010011000000: note = C1_note;
            15'b100010110100000: note = 0;
            15'b100010111000111: note = C1_note;
            15'b100011010100111: note = 0;
            15'b100011011001110: note = Ch1_note;
            15'b100011101110110: note = 0;
            15'b100011110010011: note = C1_note;
            15'b100100000111011: note = 0;
            15'b100100001011000: note = Ah_note;
            15'b100100110101000: note = 0;
            15'b100100111100010: note = Ch1_note;
            15'b100101100110010: note = 0;
            15'b100101101101100: note = Dh1_note;
            15'b100110000010100: note = 0;
            15'b100110000110001: note = F1_note;
            15'b100110110000001: note = 0;
            15'b100110110111011: note = C1_note;
            15'b100111001100011: note = 0;
            15'b100111010000000: note = Ch1_note;
            15'b100111100101000: note = 0;
            15'b100111101000101: note = C1_note;
            15'b101000010010101: note = 0;
            15'b101000011001111: note = Ch1_note;
            15'b101001000011111: note = 0;
            15'b101001001011001: note = Dh1_note;
            15'b101001100000001: note = 0;
            15'b101001100011110: note = F1_note;
            15'b101010001101110: note = 0;
            15'b101010010101000: note = Ch1_note;
            15'b101010101010000: note = 0;
            15'b101010101101101: note = C1_note;
            15'b101011000010101: note = 0;
            15'b101011000110010: note = Ch1_note;
            15'b101011110000010: note = 0;
            15'b101011110111100: note = Dh1_note;
            15'b101100001100100: note = 0;
            15'b101100010000001: note = F1_note;
            15'b101100111010001: note = 0;
            15'b101101000001011: note = C1_note;
            15'b101101010110011: note = 0;
            15'b101101011010000: note = C1_note;
            15'b101101101111000: note = 0;
            15'b101101110010101: note = C1_note;
            15'b101110011100101: note = 0;
            15'b101110100011111: note = C1_note;
            15'b101111001101111: note = 0;
            15'b101111010101001: note = C1_note;
            15'b101111101010001: note = 0;
            15'b101111101101110: note = Ch1_note;
            15'b110000000010110: note = 0;
            15'b110000000110011: note = C1_note;
            15'b110000011011011: note = 0;
            15'b110000011111000: note = Ah_note;
            15'b110000110100000: note = 0;
            15'b110000110111101: note = Ch1_note;
            15'b110001001100101: note = 0;
            15'b110001010000010: note = Ch1_note;
            15'b110001101100010: note = 0;
            15'b110001110001001: note = Ch1_note;
            15'b110010001101001: note = 0;
            15'b110010010010000: note = Ch1_note;
            15'b110010101110000: note = 0;
            15'b110010110010111: note = Ch1_note;
            15'b110011001110111: note = 0;
            15'b110011010011110: note = Ch1_note;
            15'b110011101111110: note = 0;
            15'b110011110100101: note = F1_note;
            15'b110100010000101: note = 0;
            15'b110100010101100: note = C1_note;
            15'b110100110001100: note = 0;
            15'b110100110110011: note = C1_note;
            15'b110101010010011: note = 0;
            15'b110101010111010: note = C1_note;
            15'b110101110011010: note = 0;
            15'b110101111000001: note = C1_note;
            15'b110110001101001: note = 0;
            15'b110110010000110: note = C1_note;
            15'b110110100101110: note = 0;
            15'b110110101001011: note = C1_note;
            15'b110110111110011: note = 0;
            15'b110111000010000: note = C1_note;
            15'b110111010111000: note = 0;
            15'b110111011010101: note = Ch1_note;
            15'b110111110110101: note = 0;
            15'b110111111011100: note = Ch1_note;
            15'b111000010111100: note = 0;
            15'b111000011100011: note = Ch1_note;
            15'b111000111000011: note = 0;
            15'b111000111101010: note = Ch1_note;
            15'b111001011001010: note = 0;
            15'b111001011110001: note = Ch1_note;
            15'b111001111010001: note = 0;
            15'b111001111111000: note = F1_note;
            15'b111010011011000: note = 0;
            15'b111010011111111: note = C1_note;
            15'b111010111011111: note = 0;
            15'b111011000000110: note = C1_note;
            15'b111011011100110: note = 0;
            15'b111011100001101: note = C1_note;
            15'b111011111101101: note = 0;
            15'b111100000010100: note = Ch1_note;
            15'b111100010111100: note = 0;
            15'b111100011011001: note = C1_note;
            15'b111100110000001: note = 0;
            15'b111100110011110: note = Ah_note;
            15'b111101011101110: note = 0;
            15'b111101100101000: note = Ch1_note;
            15'b111110001111000: note = 0;
            15'b111110010110010: note = Dh1_note;
            15'b111110101011010: note = 0;
            15'b111110101110111: note = F1_note;
            15'b111111011000111: note = 0;
            15'b111111100000001: note = C1_note;
            15'b111111110101001: note = 0;
            15'b111111111000110: note = Ch1_note;
            16'b1000000001101110: note = 0;
            16'b1000000010001011: note = C1_note;
            16'b1000000111011011: note = 0;
            16'b1000001000010101: note = Ch1_note;
            16'b1000001101100101: note = 0;
            16'b1000001110011111: note = Dh1_note;
            16'b1000010001000111: note = 0;
            16'b1000010001100100: note = F1_note;
            16'b1000010110110100: note = 0;
            16'b1000010111101110: note = Ch1_note;
            16'b1000011010010110: note = 0;
            16'b1000011010110011: note = C1_note;
            16'b1000011101011011: note = 0;
            16'b1000011101111000: note = Ch1_note;
            16'b1000100011001000: note = 0;
            16'b1000100100000010: note = Dh1_note;
            16'b1000100110101010: note = 0;
            16'b1000100111000111: note = F1_note;
            16'b1000101100010111: note = 0;
            16'b1000101101010001: note = C1_note;
            16'b1000101111111001: note = 0;
            16'b1000110000010110: note = C1_note;
            16'b1000110010111110: note = 0;
            16'b1000110011011011: note = C1_note;
            16'b1000111000101011: note = 0;
            16'b1000111001100101: note = C1_note;
            16'b1000111110110101: note = 0;
            16'b1000111111101111: note = C1_note;
            16'b1001000010010111: note = 0;
            16'b1001000010110100: note = Ch1_note;
            16'b1001000101011100: note = 0;
            16'b1001000101111001: note = C1_note;
            16'b1001001000100001: note = 0;
            16'b1001001000111110: note = Ah_note;
            16'b1001001110001110: note = 0;
            16'b1001001111001000: note = Gh1_note;
            16'b1001010100011000: note = 0;
            16'b1001010101010010: note = Ch1_note;
            16'b1001010111111010: note = 0;
            16'b1001011000010111: note = Ch1_note;
            16'b1001100000001111: note = 0;
            16'b1001100001100101: note = Ah_note;
            16'b1001100110110101: note = 0;
            16'b1001101010110011: note = Ch1_note;
            16'b1001101101011011: note = 0;
            16'b1001101101111000: note = Ch1_note;
            16'b1001110000100000: note = 0;
            16'b1001110000111101: note = Dh1_note;
            16'b1001110011100101: note = 0;
            16'b1001110100000010: note = F1_note;
            16'b1001110110101010: note = 0;
            16'b1001110111000111: note = Gh1_note;
            16'b1001111001101111: note = 0;
            16'b1001111010001100: note = F1_note;
            16'b1001111100110100: note = 0;
            16'b1001111101010001: note = Dh1_note;
            16'b1001111111111001: note = 0;
            16'b1010000000010110: note = Ch1_note;
            16'b1010000101100110: note = 0;
            16'b1010000110100000: note = Ch1_note;
            16'b1010001001001000: note = 0;
            16'b1010001001100101: note = Dh1_note;
            16'b1010001110110101: note = 0;
            16'b1010001111101111: note = Ch1_note;
            16'b1010010100111111: note = 0;
            16'b1010010101111001: note = F1_note;
            16'b1010011011001001: note = 0;
            16'b1010011100000011: note = Gh1_note;
            16'b1010011110101011: note = 0;
            16'b1010011111001000: note = F1_note;
            16'b1010100001110000: note = 0;
            16'b1010100010001101: note = Dh1_note;
            16'b1010100100110101: note = 0;
            16'b1010100101010010: note = Ch1_note;
            16'b1010101010100010: note = 0;
            16'b1010101011011100: note = Ah_note;
            16'b1010110000101100: note = 0;
            16'b1010110001100110: note = Gh1_note;
            16'b1010110110110110: note = 0;
            16'b1010110111110000: note = Ch1_note;
            16'b1010111010011000: note = 0;
            16'b1010111010110101: note = Ch1_note;
            16'b1011000010101101: note = 0;
            16'b1011000100000011: note = Ah_note;
            16'b1011001001010011: note = 0;
            16'b1011001101010001: note = Ch1_note;
            16'b1011001111111001: note = 0;
            16'b1011010000010110: note = Ch1_note;
            16'b1011010010111110: note = 0;
            16'b1011010011011011: note = Dh1_note;
            16'b1011010110000011: note = 0;
            16'b1011010110100000: note = F1_note;
            16'b1011011001001000: note = 0;
            16'b1011011001100101: note = Gh1_note;
            16'b1011011100001101: note = 0;
            16'b1011011100101010: note = F1_note;
            16'b1011011111010010: note = 0;
            16'b1011011111101111: note = Dh1_note;
            16'b1011100010010111: note = 0;
            16'b1011100010110100: note = Ch1_note;
            16'b1011101000000100: note = 0;
            16'b1011101000111110: note = Ch1_note;
            16'b1011101011100110: note = 0;
            16'b1011101100000011: note = Dh1_note;
            16'b1011110001010011: note = 0;
            16'b1011110010001101: note = Ch1_note;
            16'b1011110111011101: note = 0;
            16'b1011111000010111: note = F1_note;
            16'b1011111101100111: note = 0;
            16'b1011111110100001: note = Gh1_note;
            16'b1100000001001001: note = 0;
            16'b1100000001100110: note = F1_note;
            16'b1100000100001110: note = 0;
            16'b1100000100101011: note = Dh1_note;
            16'b1100000111010011: note = 0;
            16'b1100000111110000: note = Ch1_note;
            16'b1100001101000000: note = 0;
            16'b1100001101111010: note = Ah_note;
            16'b1100010000100010: note = 0;
            16'b1100010000111111: note = Ah_note;
            16'b1100010011100111: note = 0;
            16'b1100010100000100: note = Ch1_note;
            16'b1100010101110011: note = 0;
            16'b1100010110000111: note = Ch1_note;
            16'b1100010111110110: note = 0;
            16'b1100011000001010: note = Ch1_note;
            16'b1100011001111001: note = 0;
            16'b1100011010001101: note = Ch1_note;
            16'b1100011011111100: note = 0;
            16'b1100011100010000: note = Ch1_note;
            16'b1100011101111111: note = 0;
            16'b1100011110010011: note = Ch1_note;
            16'b1100100000000010: note = 0;
            16'b1100100000010110: note = Dh1_note;
            16'b1100100101100110: note = 0;
            16'b1100100110100000: note = F1_note;
            16'b1100101000001111: note = 0;
            16'b1100101000100011: note = C1_note;
            16'b1100101010010010: note = 0;
            16'b1100101010100110: note = C1_note;
            16'b1100101100010101: note = 0;
            16'b1100101100101001: note = C1_note;
            16'b1100101110011000: note = 0;
            16'b1100101110101100: note = C1_note;
            16'b1100110000011011: note = 0;
            16'b1100110000101111: note = C1_note;
            16'b1100110010011110: note = 0;
            16'b1100110010110010: note = Ch1_note;
            16'b1100111000000010: note = 0;
            16'b1100111000111100: note = F1_note;
            16'b1100111100111000: note = 0;
            16'b1100111101100100: note = C1_note;
            16'b1101000000101000: note = 0;
            16'b1101000001001001: note = C1_note;
            16'b1101000010111000: note = 0;
            16'b1101000011001100: note = C1_note;
            16'b1101000100111011: note = 0;
            16'b1101000101001111: note = Ch1_note;
            16'b1101001010011111: note = 0;
            16'b1101001011011001: note = F1_note;
            16'b1101001101001000: note = 0;
            16'b1101001101011100: note = F1_note;
            16'b1101001111001011: note = 0;
            16'b1101001111011111: note = F1_note;
            16'b1101010001001110: note = 0;
            16'b1101010001100010: note = C1_note;
            16'b1101010110110010: note = 0;
            16'b1101010111101100: note = Dh1_note;
            16'b1101011100111100: note = 0;
            16'b1101011101110110: note = Ch1_note;
            16'b1101100011000110: note = 0;
            16'b1101100100000000: note = F1_note;
            16'b1101100101101111: note = 0;
            16'b1101100110000011: note = F1_note;
            16'b1101100111110010: note = 0;
            16'b1101101000000110: note = Dh1_note;
            16'b1101101001110101: note = 0;
            16'b1101101010001001: note = Ch1_note;
            16'b1101101011111000: note = 0;
            16'b1101101100001100: note = C1_note;
            16'b1101101101111011: note = 0;
            16'b1101101110001111: note = C1_note;
            16'b1101101111111110: note = 0;
            16'b1101110000010010: note = Dh1_note;
            16'b1101110101100010: note = 0;
            16'b1101110110011100: note = Ch1_note;
            16'b1101111011101100: note = 0;
            16'b1101111100100110: note = F1_note;
            16'b1110000001110110: note = 0;
            16'b1110000010110000: note = C1_note;
            16'b1110000100011111: note = 0;
            16'b1110000100110011: note = C1_note;
            16'b1110000110100010: note = 0;
            16'b1110000110110110: note = C1_note;
            16'b1110001000100101: note = 0;
            16'b1110001000111001: note = Dh1_note;
            16'b1110001110001001: note = 0;
            16'b1110001111000011: note = Ch1_note;
            16'b1110010100010011: note = 0;
            16'b1110010101001101: note = F1_note;
            16'b1110010111110101: note = 0;
            16'b1110011000010010: note = F1_note;
            16'b1110011010111010: note = 0;
            16'b1110011011010111: note = C1_note;
            16'b1110011101000110: note = 0;
            16'b1110011101011010: note = C1_note;
            16'b1110011111001001: note = 0;
            16'b1110011111011101: note = C1_note;
            16'b1110100001001100: note = 0;
            16'b1110100001100000: note = Dh1_note;
            16'b1110100110110000: note = 0;
            16'b1110100111101010: note = Ch1_note;
            16'b1110101100111010: note = 0;
            16'b1110101101110100: note = F1_note;
            16'b1110110000011100: note = 0;
            16'b1110110000111001: note = C1_note;
            16'b1110110011100001: note = 0;
            16'b1110110011111110: note = C1_note;
            16'b1110110101101101: note = 0;
            16'b1110110110000001: note = C1_note;
            16'b1110110111110000: note = 0;
            16'b1110111000000100: note = C1_note;
            16'b1110111001110011: note = 0;
            16'b1110111010000111: note = Dh1_note;
            16'b1110111111010111: note = 0;
            16'b1111000000010001: note = Ch1_note;
            16'b1111000101100001: note = 0;
            16'b1111000110011011: note = F1_note;
            16'b1111001001000011: note = 0;
            16'b1111001001100000: note = C1_note;
            16'b1111001100001000: note = 0;
            16'b1111001100100101: note = C1_note;
            16'b1111001110010100: note = 0;
            16'b1111001110101000: note = C1_note;
            16'b1111010000010111: note = 0;
            16'b1111010000101011: note = C1_note;
            16'b1111010010011010: note = 0;
            16'b1111010010101110: note = C1_note;
            16'b1111010111111110: note = 0;
            16'b1111011000111000: note = Ah_note;
            16'b1111100000110000: note = 0;
            16'b1111100010000110: note = Ch1_note;
            16'b1111100100101110: note = 0;
            16'b1111100101001011: note = Ch1_note;
            16'b1111100111110011: note = 0;
            16'b1111101000010000: note = Dh1_note;
            16'b1111101010111000: note = 0;
            16'b1111101011010101: note = Ch1_note;
            16'b1111101101111101: note = 0;
            16'b1111101110011010: note = Dh1_note;
            16'b1111110011101010: note = 0;
            16'b1111110100100100: note = C1_note;
            16'b1111110111001100: note = 0;
            16'b1111110111101001: note = C1_note;
            16'b1111111010010001: note = 0;
            16'b1111111010101110: note = C1_note;
            16'b1111111101010110: note = 0;
            16'b1111111101110011: note = C1_note;
            17'b10000000000011011: note = 0;
            17'b10000000000111000: note = C1_note;
            17'b10000000011100000: note = 0;
            17'b10000000011111101: note = Ch1_note;
            17'b10000001001001101: note = 0;
            17'b10000001010000111: note = Ch1_note;
            17'b10000001100101111: note = 0;
            17'b10000001101001100: note = Ch1_note;
            17'b10000001111110100: note = 0;
            17'b10000010000010001: note = Ch1_note;
            17'b10000010010111001: note = 0;
            17'b10000010011010110: note = Ch1_note;
            17'b10000010101111110: note = 0;
            17'b10000010110011011: note = Ch1_note;
            17'b10000011001000011: note = 0;
            17'b10000011001100000: note = Dh1_note;
            17'b10000011100001000: note = 0;
            17'b10000011100100101: note = Ch1_note;
            17'b10000011111001101: note = 0;
            17'b10000011111101010: note = Dh1_note;
            17'b10000100100111010: note = 0;
            17'b10000100101110100: note = C1_note;
            17'b10000101000011100: note = 0;
            17'b10000101000111001: note = C1_note;
            17'b10000101011100001: note = 0;
            17'b10000101011111110: note = C1_note;
            17'b10000101110100110: note = 0;
            17'b10000101111000011: note = C1_note;
            17'b10000110001101011: note = 0;
            17'b10000110010001000: note = C1_note;
            17'b10000110100110000: note = 0;
            17'b10000110101001101: note = Ch1_note;
            17'b10000111010011101: note = 0;
            17'b10000111011010111: note = Ch2_note;
            17'b10000111101111111: note = 0;
            17'b10000111110011100: note = Ch2_note;
            17'b10001000001000100: note = 0;
            17'b10001000001100001: note = Ch2_note;
            17'b10001000100001001: note = 0;
            17'b10001000100100110: note = Ch2_note;
            17'b10001000111001110: note = 0;
            17'b10001000111101011: note = Ch2_note;
            17'b10001001010010011: note = 0;
            17'b10001001010110000: note = Dh2_note;
            17'b10001001101011000: note = 0;
            17'b10001001101110101: note = Ch2_note;
            17'b10001010000011101: note = 0;
            17'b10001010000111010: note = Dh2_note;
            17'b10001010110001010: note = 0;
            17'b10001010111000100: note = C2_note;
            17'b10001011001101100: note = 0;
            17'b10001011010001001: note = C2_note;
            17'b10001011100110001: note = 0;
            17'b10001011101001110: note = C2_note;
            17'b10001011111110110: note = 0;
            17'b10001100000010011: note = C2_note;
            17'b10001100010111011: note = 0;
            17'b10001100011011000: note = C2_note;
            17'b10001100110000000: note = 0;
            17'b10001100110011101: note = Ch2_note;
            17'b10001101011101101: note = 0;
            17'b10001101100100111: note = Ch2_note;
            17'b10001101111001111: note = 0;
            17'b10001101111101100: note = Ch2_note;
            17'b10001110010010100: note = 0;
            17'b10001110010110001: note = Ch2_note;
            17'b10001110101011001: note = 0;
            17'b10001110101110110: note = Ch2_note;
            17'b10001111000011110: note = 0;
            17'b10001111000111011: note = Ch2_note;
            17'b10001111011100011: note = 0;
            17'b10001111100000000: note = Dh2_note;
            17'b10001111110101000: note = 0;
            17'b10001111111000101: note = Ch2_note;
            17'b10010000001101101: note = 0;
            17'b10010000010001010: note = Dh2_note;
            17'b10010000111011010: note = 0;
            17'b10010001000010100: note = C2_note;
            17'b10010001010111100: note = 0;
            17'b10010001011011001: note = C2_note;
            17'b10010001110000001: note = 0;
            17'b10010001110011110: note = C2_note;
            17'b10010010001000110: note = 0;
            17'b10010010001100011: note = C2_note;
            17'b10010010100001011: note = 0;
            17'b10010010100101000: note = C2_note;
            17'b10010010111010000: note = 0;
            17'b10010010111101101: note = Ch2_note;
            17'b10010011100111101: note = 0;
            17'b10010011101110111: note = Ch1_note;
            17'b10010100001010111: note = 0;
            17'b10010100001111110: note = Ch1_note;
            17'b10010100101011110: note = 0;
            17'b10010100110000101: note = Ch1_note;
            17'b10010101001100101: note = 0;
            17'b10010101010001100: note = Ch1_note;
            17'b10010101101101100: note = 0;
            17'b10010101110010011: note = Ch1_note;
            17'b10010110001110011: note = 0;
            17'b10010110010011010: note = F1_note;
            17'b10010110101111010: note = 0;
            17'b10010110110100001: note = C1_note;
            17'b10010111010000001: note = 0;
            17'b10010111010101000: note = C1_note;
            17'b10010111110001000: note = 0;
            17'b10010111110101111: note = C1_note;
            17'b10011000010001111: note = 0;
            17'b10011000010110110: note = C1_note;
            17'b10011000101011110: note = 0;
            17'b10011000101111011: note = C1_note;
            17'b10011001000100011: note = 0;
            17'b10011001001000000: note = C1_note;
            17'b10011001011101000: note = 0;
            17'b10011001100000101: note = C1_note;
            17'b10011001110101101: note = 0;
            17'b10011001111001010: note = Ch1_note;
            17'b10011010010101010: note = 0;
            17'b10011010011010001: note = Ch1_note;
            17'b10011010110110001: note = 0;
            17'b10011010111011000: note = Ch1_note;
            17'b10011011010111000: note = 0;
            17'b10011011011011111: note = Ch1_note;
            17'b10011011110111111: note = 0;
            17'b10011011111100110: note = Ch1_note;
            17'b10011100011000110: note = 0;
            17'b10011100011101101: note = F1_note;
            17'b10011100111001101: note = 0;
            17'b10011100111110100: note = C1_note;
            17'b10011101011010100: note = 0;
            17'b10011101011111011: note = C1_note;
            17'b10011101111011011: note = 0;
            17'b10011110000000010: note = C1_note;
            17'b10011110011100010: note = 0;
            17'b10011110100001001: note = Ch1_note;
            17'b10011110110110001: note = 0;
            17'b10011110111001110: note = C1_note;
            17'b10011111001110110: note = 0;
            17'b10011111010010011: note = Ah_note;
            17'b10011111111100011: note = 0;
            17'b10100000000011101: note = Ch1_note;
            17'b10100000101101101: note = 0;
            17'b10100000110100111: note = Dh1_note;
            17'b10100001001001111: note = 0;
            17'b10100001001101100: note = F1_note;
            17'b10100001110111100: note = 0;
            17'b10100001111110110: note = C1_note;
            17'b10100010010011110: note = 0;
            17'b10100010010111011: note = Ch1_note;
            17'b10100010101100011: note = 0;
            17'b10100010110000000: note = C1_note;
            17'b10100011011010000: note = 0;
            17'b10100011100001010: note = Ch1_note;
            17'b10100100001011010: note = 0;
            17'b10100100010010100: note = Dh1_note;
            17'b10100100100111100: note = 0;
            17'b10100100101011001: note = F1_note;
            17'b10100101010101001: note = 0;
            17'b10100101011100011: note = Ch1_note;
            17'b10100101110001011: note = 0;
            17'b10100101110101000: note = C1_note;
            17'b10100110001010000: note = 0;
            17'b10100110001101101: note = Ch1_note;
            17'b10100110110111101: note = 0;
            17'b10100110111110111: note = Dh1_note;
            17'b10100111010011111: note = 0;
            17'b10100111010111100: note = F1_note;
            17'b10101000000001100: note = 0;
            17'b10101000001000110: note = C1_note;
            17'b10101000011101110: note = 0;
            17'b10101000100001011: note = C1_note;
            17'b10101000110110011: note = 0;
            17'b10101000111010000: note = C1_note;
            17'b10101001100100000: note = 0;
            17'b10101001101011010: note = C1_note;
            17'b10101010010101010: note = 0;
            17'b10101010011100100: note = C1_note;
            17'b10101010110001100: note = 0;
            17'b10101010110101001: note = Ch1_note;
            17'b10101011001010001: note = 0;
            17'b10101011001101110: note = C1_note;
            17'b10101011100010110: note = 0;
            17'b10101011100110011: note = Ah_note;
            17'b10101011111011011: note = 0;
            17'b10101011111111000: note = Ch1_note;
            17'b10101100010100000: note = 0;
            17'b10101100010111101: note = Ch1_note;
            17'b10101100110011101: note = 0;
            17'b10101100111000100: note = Ch1_note;
            17'b10101101010100100: note = 0;
            17'b10101101011001011: note = Ch1_note;
            17'b10101101110101011: note = 0;
            17'b10101101111010010: note = Ch1_note;
            17'b10101110010110010: note = 0;
            17'b10101110011011001: note = Ch1_note;
            17'b10101110110111001: note = 0;
            17'b10101110111100000: note = F1_note;
            17'b10101111011000000: note = 0;
            17'b10101111011100111: note = C1_note;
            17'b10101111111000111: note = 0;
            17'b10101111111101110: note = C1_note;
            17'b10110000011001110: note = 0;
            17'b10110000011110101: note = C1_note;
            17'b10110000111010101: note = 0;
            17'b10110000111111100: note = C1_note;
            17'b10110001010100100: note = 0;
            17'b10110001011000001: note = C1_note;
            17'b10110001101101001: note = 0;
            17'b10110001110000110: note = C1_note;
            17'b10110010000101110: note = 0;
            17'b10110010001001011: note = C1_note;
            17'b10110010011110011: note = 0;
            17'b10110010100010000: note = Ch1_note;
            17'b10110010111110000: note = 0;
            17'b10110011000010111: note = Ch1_note;
            17'b10110011011110111: note = 0;
            17'b10110011100011110: note = Ch1_note;
            17'b10110011111111110: note = 0;
            17'b10110100000100101: note = Ch1_note;
            17'b10110100100000101: note = 0;
            17'b10110100100101100: note = Ch1_note;
            17'b10110101000001100: note = 0;
            17'b10110101000110011: note = F1_note;
            17'b10110101100010011: note = 0;
            17'b10110101100111010: note = C1_note;
            17'b10110110000011010: note = 0;
            17'b10110110001000001: note = C1_note;
            17'b10110110100100001: note = 0;
            17'b10110110101001000: note = C1_note;
            17'b10110111000101000: note = 0;
            17'b10110111001001111: note = Ch1_note;
            17'b10110111011110111: note = 0;
            17'b10110111100010100: note = C1_note;
            17'b10110111110111100: note = 0;
            17'b10110111111011001: note = Ah_note;
            17'b10111000100101001: note = 0;
            17'b10111000101100011: note = Ch1_note;
            17'b10111001010110011: note = 0;
            17'b10111001011101101: note = Dh1_note;
            17'b10111001110010101: note = 0;
            17'b10111001110110010: note = F1_note;
            17'b10111010100000010: note = 0;
            17'b10111010100111100: note = C1_note;
            17'b10111010111100100: note = 0;
            17'b10111011000000001: note = Ch1_note;
            17'b10111011010101001: note = 0;
            17'b10111011011000110: note = C1_note;
            17'b10111100000010110: note = 0;
            17'b10111100001010000: note = Ch1_note;
            17'b10111100110100000: note = 0;
            17'b10111100111011010: note = Dh1_note;
            17'b10111101010000010: note = 0;
            17'b10111101010011111: note = F1_note;
            17'b10111101111101111: note = 0;
            17'b10111110000101001: note = Ch1_note;
            17'b10111110011010001: note = 0;
            17'b10111110011101110: note = C1_note;
            17'b10111110110010110: note = 0;
            17'b10111110110110011: note = Ch1_note;
            17'b10111111100000011: note = 0;
            17'b10111111100111101: note = Dh1_note;
            17'b10111111111100101: note = 0;
            17'b11000000000000010: note = F1_note;
            17'b11000000101010010: note = 0;
            17'b11000000110001100: note = C1_note;
            17'b11000001000110100: note = 0;
            17'b11000001001010001: note = C1_note;
            17'b11000001011111001: note = 0;
            17'b11000001100010110: note = C1_note;
            17'b11000010001100110: note = 0;
            17'b11000010010100000: note = C1_note;
            17'b11000010111110000: note = 0;
            17'b11000011000101010: note = C1_note;
            17'b11000011011010010: note = 0;
            17'b11000011011101111: note = Ch1_note;
            17'b11000011110010111: note = 0;
            17'b11000011110110100: note = C1_note;
            17'b11000100001011100: note = 0;
            17'b11000100001111001: note = Ah_note;
            17'b11000100100100001: note = 0;
            17'b11000100100111110: note = Fh1_note;
            17'b11000100111100110: note = 0;
            17'b11000101000000011: note = F1_note;
            17'b11000110101001100: note = 0;
            17'b11000110111011011: note = Ch1_note;
            17'b11000111010000011: note = 0;
            17'b11000111010100000: note = Dh1_note;
            17'b11000111111110000: note = 0;
            17'b11001000000101010: note = Ch1_note;
            17'b11001001011001010: note = 0;
            17'b11001001100111101: note = F1_note;
            17'b11001001111100101: note = 0;
            17'b11001010000000010: note = Fh1_note;
            17'b11001010010101010: note = 0;
            17'b11001010011000111: note = F1_note;
            17'b11001010101101111: note = 0;
            17'b11001010110001100: note = Dh1_note;
            17'b11001011000110100: note = 0;
            17'b11001011001010001: note = F1_note;
            17'b11001100110011010: note = 0;
            17'b11001101000101001: note = Ch1_note;
            17'b11001101011010001: note = 0;
            17'b11001101011101110: note = Dh1_note;
            17'b11001101110010110: note = 0;
            17'b11001101110110011: note = Ch1_note;
            17'b11001110100000011: note = 0;
            17'b11001110100111101: note = Dh1_note;
            17'b11001111010001101: note = 0;
            17'b11001111011000111: note = F1_note;
            17'b11001111101101111: note = 0;
            17'b11001111110001100: note = F1_note;
            17'b11010000000110100: note = 0;
            17'b11010000001010001: note = Dh1_note;
            17'b11010000011111001: note = 0;
            17'b11010000100010110: note = F1_note;
            17'b11010000110111110: note = 0;
            17'b11010000111011011: note = Dh1_note;
            17'b11010001010000011: note = 0;
            17'b11010001010100000: note = F1_note;
            17'b11010010111101001: note = 0;
            17'b11010011001111000: note = Ch1_note;
            17'b11010011100100000: note = 0;
            17'b11010011100111101: note = Dh1_note;
            17'b11010100010001101: note = 0;
            17'b11010100011000111: note = Ch1_note;
            17'b11010101010111111: note = 0;
            17'b11010101100010101: note = Dh1_note;
            17'b11010101110111101: note = 0;
            17'b11010101111011010: note = F1_note;
            17'b11010110010000010: note = 0;
            17'b11010110010011111: note = F1_note;
            17'b11010110101000111: note = 0;
            17'b11010110101100100: note = F1_note;
            17'b11010111000001100: note = 0;
            17'b11010111000101001: note = Dh1_note;
            17'b11010111011010001: note = 0;
            17'b11010111011101110: note = F1_note;
            17'b11011000000111110: note = 0;
            17'b11011000001111000: note = Ch1_note;
            17'b11011001001110000: note = 0;
            17'b11011001011000110: note = Ch1_note;
            17'b11011001101101110: note = 0;
            17'b11011001110001011: note = Dh1_note;
            17'b11011010000110011: note = 0;
            17'b11011010001010000: note = Ch1_note;
            17'b11011010110100000: note = 0;
            17'b11011010111011010: note = Ah_note;
            17'b11011100100100011: note = 0;
            17'b11011100110110010: note = F1_note;
            17'b11011101100000010: note = 0;
            17'b11011101100111100: note = F1_note;
            17'b11011101111100100: note = 0;
            17'b11011110000000001: note = Ch1_note;
            17'b11011110010101001: note = 0;
            17'b11011110011000110: note = Dh1_note;
            17'b11011111000010110: note = 0;
            17'b11011111001010000: note = Ah1_note;
            17'b11011111011111000: note = 0;
            17'b11011111100010101: note = Ch2_note;
            17'b11011111110111101: note = 0;
            17'b11011111111011010: note = Ch2_note;
            17'b11100000100101010: note = 0;
            17'b11100000101100100: note = Ah1_note;
            17'b11100001010110100: note = 0;
            17'b11100001011101110: note = Ch2_note;
            17'b11100010000111110: note = 0;
            17'b11100010001111000: note = Ah1_note;
            17'b11100010100100000: note = 0;
            17'b11100010100111101: note = Ch2_note;
            17'b11100010111100101: note = 0;
            17'b11100011000000010: note = Ch2_note;
            17'b11100011101010010: note = 0;
            17'b11100011110001100: note = Ah1_note;
            17'b11100100011011100: note = 0;
            17'b11100100100010110: note = Ch2_note;
            17'b11100101001100110: note = 0;
            17'b11100101010100000: note = Ah1_note;
            17'b11100101101001000: note = 0;
            17'b11100101101100101: note = Ch2_note;
            17'b11100110000001101: note = 0;
            17'b11100110000101010: note = Ch2_note;
            17'b11100110101111010: note = 0;
            17'b11100110110110100: note = Ah1_note;
            17'b11100111001011100: note = 0;
            17'b11100111001111001: note = Ch2_note;
            17'b11100111100100001: note = 0;
            17'b11100111100111110: note = Ch2_note;
            17'b11101000010001110: note = 0;
            17'b11101000011001000: note = F1_note;
            17'b11101000101110000: note = 0;
            17'b11101000110001101: note = Fh1_note;
            17'b11101001000110101: note = 0;
            17'b11101001001010010: note = F1_note;
            17'b11101001011111010: note = 0;
            17'b11101001100010111: note = Dh1_note;
            17'b11101001110111111: note = 0;
            17'b11101001111011100: note = F1_note;
            17'b11101010010000100: note = 0;
            17'b11101010010100001: note = Ch1_note;
            17'b11101010101001001: note = 0;
            17'b11101010101100110: note = Dh1_note;
            17'b11101100101010111: note = 0;
            17'b11101101000000011: note = Ch2_note;
            17'b11101101010101011: note = 0;
            17'b11101101011001000: note = Dh2_note;
            17'b11101101101110000: note = 0;
            17'b11101101110001101: note = C2_note;
            17'b11101110011011101: note = 0;
            17'b11101110100010111: note = F2_note;
            17'b11101110110111111: note = 0;
            17'b11101110111011100: note = Fh2_note;
            17'b11101111010000100: note = 0;
            17'b11101111010100001: note = F2_note;
            17'b11101111101001001: note = 0;
            17'b11101111101100110: note = Dh2_note;
            17'b11110000000001110: note = 0;
            17'b11110000000101011: note = F2_note;
            17'b11110000011010011: note = 0;
            17'b11110000011110000: note = Ch2_note;
            17'b11110000110011000: note = 0;
            17'b11110000110110101: note = Dh2_note;
            17'b11110010001010101: note = 0;
            17'b11110010011001000: note = Ch2_note;
            17'b11110011000011000: note = 0;
            17'b11110011001010010: note = Ch2_note;
            17'b11110011011111010: note = 0;
            17'b11110011100010111: note = Dh2_note;
            17'b11110011110111111: note = 0;
            17'b11110011111011100: note = C2_note;
            17'b11110100100101100: note = 0;
            17'b11110100101100110: note = C2_note;
            17'b11110101000001110: note = 0;
            17'b11110101000101011: note = Dh2_note;
            17'b11110101011010011: note = 0;
            17'b11110101011110000: note = F2_note;
            17'b11110110001000000: note = 0;
        endcase
    end   
    //my_war
    else if (sw_state == 4'b0011) begin
        case (counter_sec) 
            2'b11: note = Dh1_note;
            10'b1001001001: note = 0;
            10'b1010101101: note = E1_note;
            11'b10011110110: note = 0;
            11'b10101011010: note = Dh1_note;
            11'b11110100011: note = 0;
            12'b100000000111: note = C2_note;
            12'b100100101011: note = 0;
            12'b100101011110: note = Gh2_note;
            12'b101010000010: note = 0;
            12'b101010110101: note = Dh1_note;
            12'b110011111110: note = 0;
            12'b110101100010: note = E1_note;
            12'b111110101011: note = 0;
            13'b1000000001111: note = Dh1_note;
            13'b1001001011000: note = 0;
            13'b1001010111100: note = Ch3_note;
            13'b1001100000101: note = 0;
            13'b1001100010010: note = Ch2_note;
            13'b1001101011011: note = 0;
            13'b1001101101000: note = B2_note;
            13'b1001110110001: note = 0;
            13'b1001110111110: note = B1_note;
            13'b1010000000111: note = 0;
            13'b1010000010100: note = A2_note;
            13'b1010001011101: note = 0;
            13'b1010001101010: note = A1_note;
            13'b1010010110011: note = 0;
            13'b1010011000000: note = Gh2_note;
            13'b1010100001001: note = 0;
            13'b1010100010110: note = Gh1_note;
            13'b1010101011111: note = 0;
            13'b1010101100111: note = Ch1_note;
            13'b1011010011011: note = 0;
            13'b1011010111101: note = E1_note;
            13'b1011111010010: note = 0;
            13'b1100000010100: note = E1_note;
            13'b1100010100110: note = 0;
            13'b1100010111111: note = Ch1_note;
            13'b1100111100011: note = 0;
            13'b1101000010110: note = Ch1_note;
            13'b1101010101000: note = 0;
            13'b1101011000001: note = Ch1_note;
            13'b1101101010011: note = 0;
            13'b1101101101100: note = Gh1_note;
            13'b1101111111110: note = 0;
            13'b1110000010111: note = Gh1_note;
            13'b1110010101001: note = 0;
            13'b1110011000010: note = Gh1_note;
            13'b1110101010100: note = 0;
            13'b1110101101101: note = Gh1_note;
            13'b1111010010001: note = 0;
            13'b1111011000100: note = E1_note;
            13'b1111101010110: note = 0;
            13'b1111101101111: note = Dh1_note;
            14'b10000000000001: note = 0;
            14'b10000000011010: note = Ch1_note;
            14'b10001001100011: note = 0;
            14'b10001011000111: note = E1_note;
            14'b10001101011001: note = 0;
            14'b10001101110010: note = Ch1_note;
            14'b10010010010110: note = 0;
            14'b10010011001001: note = Ch1_note;
            14'b10010101011011: note = 0;
            14'b10010101110100: note = Ch1_note;
            14'b10011000000110: note = 0;
            14'b10011000011111: note = Gh1_note;
            14'b10011010110001: note = 0;
            14'b10011011001010: note = Gh1_note;
            14'b10011101011100: note = 0;
            14'b10011101110101: note = Gh1_note;
            14'b10100000000111: note = 0;
            14'b10100000100000: note = Ch2_note;
            14'b10100010110010: note = 0;
            14'b10100011001011: note = B1_note;
            14'b10100101011101: note = 0;
            14'b10100101110110: note = A1_note;
            14'b10101000001000: note = 0;
            14'b10101000100001: note = Gh1_note;
            14'b10101010110011: note = 0;
            14'b10101011001100: note = Ch1_note;
            14'b10110000000000: note = 0;
            14'b10110000100010: note = E1_note;
            14'b10110100110111: note = 0;
            14'b10110101111001: note = E1_note;
            14'b10111000001011: note = 0;
            14'b10111000100100: note = Ch1_note;
            14'b10111101001000: note = 0;
            14'b10111101111011: note = Ch1_note;
            14'b11000000001101: note = 0;
            14'b11000000100110: note = Ch1_note;
            14'b11000010111000: note = 0;
            14'b11000011010001: note = Gh1_note;
            14'b11000101100011: note = 0;
            14'b11000101111100: note = Gh1_note;
            14'b11001000001110: note = 0;
            14'b11001000100111: note = Gh1_note;
            14'b11001010111001: note = 0;
            14'b11001011010010: note = Gh1_note;
            14'b11001111110110: note = 0;
            14'b11010000101001: note = E1_note;
            14'b11010010111011: note = 0;
            14'b11010011010100: note = Dh1_note;
            14'b11010101100110: note = 0;
            14'b11010101111111: note = Ch1_note;
            14'b11011010100011: note = 0;
            14'b11011011010110: note = Ch2_note;
            14'b11100000001010: note = 0;
            14'b11100000101101: note = Ch1_note;
            14'b11100101010001: note = 0;
            14'b11100110000100: note = Ch2_note;
            14'b11101010111000: note = 0;
            14'b11101011011011: note = Ch1_note;
            14'b11101101101101: note = 0;
            14'b11101110000110: note = Ch2_note;
            14'b11110000011000: note = 0;
            14'b11110000110001: note = Ch2_note;
            14'b11110011000011: note = 0;
            14'b11110011011100: note = Ch2_note;
            14'b11110101101110: note = 0;
            14'b11110110000111: note = Ch2_note;
            14'b11111000011001: note = 0;
            14'b11111000110010: note = B1_note;
            14'b11111011000100: note = 0;
            14'b11111011011101: note = A1_note;
            14'b11111101101111: note = 0;
            14'b11111110001000: note = Ch2_note;
            14'b11111111010001: note = 0;
            14'b11111111011110: note = Dh2_note;
            15'b100000000100111: note = 0;
            15'b100000000110100: note = E2_note;
            15'b100000011000110: note = 0;
            15'b100000011011111: note = Dh2_note;
            15'b100000101110001: note = 0;
            15'b100000110001010: note = Fh2_note;
            15'b100001000011100: note = 0;
            15'b100001000110101: note = E2_note;
            15'b100001011000111: note = 0;
            15'b100001011100000: note = Gh2_note;
            15'b100001101110010: note = 0;
            15'b100001110001011: note = Fh2_note;
            15'b100010000011101: note = 0;
            15'b100010000110110: note = A2_note;
            15'b100010011001000: note = 0;
            15'b100010011100001: note = Gh2_note;
            15'b100010101110011: note = 0;
            15'b100010110001100: note = Fh2_note;
            15'b100011000011110: note = 0;
            15'b100011000110111: note = Gh2_note;
            15'b100011011001001: note = 0;
            15'b100011011100010: note = E2_note;
            15'b100011101110100: note = 0;
            15'b100011110001101: note = Dh2_note;
            15'b100100000011111: note = 0;
            15'b100100000111000: note = E2_note;
            15'b100100011001010: note = 0;
            15'b100100011100011: note = Gh2_note;
            15'b100100101110101: note = 0;
            15'b100100110001110: note = Dh2_note;
            15'b100101000100000: note = 0;
            15'b100101000111001: note = Gh2_note;
            15'b100101011001011: note = 0;
            15'b100101011100100: note = Ch2_note;
            15'b100101101110110: note = 0;
            15'b100101110001111: note = Gh1_note;
            15'b100110000100001: note = 0;
            15'b100110000111010: note = Ch2_note;
            15'b100110011001100: note = 0;
            15'b100110011100101: note = Dh2_note;
            15'b100110101110111: note = 0;
            15'b100110110010000: note = E2_note;
            15'b100111000100010: note = 0;
            15'b100111000111011: note = Gh1_note;
            15'b100111011001101: note = 0;
            15'b100111011100110: note = Dh2_note;
            15'b100111101111000: note = 0;
            15'b100111110010001: note = Gh1_note;
            15'b101000000100011: note = 0;
            15'b101000000111100: note = Ch2_note;
            15'b101000011001110: note = 0;
            15'b101000011100111: note = Gh1_note;
            15'b101000101111001: note = 0;
            15'b101000110010010: note = Ch2_note;
            15'b101001000100100: note = 0;
            15'b101001000111101: note = Gh1_note;
            15'b101001011001111: note = 0;
            15'b101001011101000: note = Ch2_note;
            15'b101001101111010: note = 0;
            15'b101001110010011: note = B1_note;
            15'b101010000100101: note = 0;
            15'b101010000111110: note = Gh2_note;
            15'b101010101100010: note = 0;
            15'b101010110010101: note = E3_note;
            15'b101011010111001: note = 0;
            15'b101011011101100: note = Fh3_note;
            15'b101011101111110: note = 0;
            15'b101011110010111: note = Dh3_note;
            15'b101100010111011: note = 0;
            15'b101100011101110: note = E3_note;
            15'b101101000010010: note = 0;
            15'b101101001000101: note = Ch3_note;
            15'b101101101101001: note = 0;
            15'b101101110011100: note = Dh3_note;
            15'b101110011000000: note = 0;
            15'b101110011110011: note = A2_note;
            15'b101111000010111: note = 0;
            15'b101111001001010: note = Gh2_note;
            15'b101111101101110: note = 0;
            15'b101111110100001: note = Gh2_note;
            15'b110000000110011: note = 0;
            15'b110000001001100: note = E3_note;
            15'b110000101110000: note = 0;
            15'b110000110100011: note = Fh3_note;
            15'b110001000110101: note = 0;
            15'b110001001001110: note = Dh3_note;
            15'b110001101110010: note = 0;
            15'b110001110100101: note = E3_note;
            15'b110010011001001: note = 0;
            15'b110010011111100: note = Ch3_note;
            15'b110011000100000: note = 0;
            15'b110011001010011: note = B3_note;
            15'b110011101110111: note = 0;
            15'b110011110101010: note = Ch4_note;
            15'b110100101100001: note = 0;
            15'b110100110101011: note = Gh2_note;
            15'b110101011001111: note = 0;
            15'b110101100000010: note = E3_note;
            15'b110110000100110: note = 0;
            15'b110110001011001: note = Fh3_note;
            15'b110110011101011: note = 0;
            15'b110110100000100: note = Dh3_note;
            15'b110111000101000: note = 0;
            15'b110111001011011: note = E3_note;
            15'b110111101111111: note = 0;
            15'b110111110110010: note = Ch3_note;
            15'b111000011010110: note = 0;
            15'b111000100001001: note = Dh3_note;
            15'b111001000101101: note = 0;
            15'b111001001100000: note = A2_note;
            15'b111001110000100: note = 0;
            15'b111001110110111: note = Gh2_note;
            15'b111010101101110: note = 0;
            15'b111010110111000: note = E2_note;
            15'b111011011011100: note = 0;
            15'b111011100001111: note = Gh2_note;
            15'b111011110100001: note = 0;
            15'b111011110111010: note = Dh2_note;
            15'b111100011011110: note = 0;
            15'b111100100010001: note = Gh2_note;
            15'b111101000110101: note = 0;
            15'b111101001101000: note = E1_note;
            15'b111101011111010: note = 0;
            15'b111110110110111: note = D3_note;
            15'b111111000000000: note = 0;
            15'b111111000001101: note = D2_note;
            15'b111111001010110: note = 0;
            15'b111111001100011: note = C3_note;
            15'b111111010101100: note = 0;
            15'b111111010111001: note = C2_note;
            15'b111111100000010: note = 0;
            15'b111111100001111: note = Ah2_note;
            15'b111111101011000: note = 0;
            15'b111111101100101: note = Ah1_note;
            15'b111111110101110: note = 0;
            15'b111111110111011: note = A2_note;
            16'b1000000000000100: note = 0;
            16'b1000000000010001: note = A1_note;
            16'b1000000001011010: note = 0;
            16'b1000000001100111: note = D1_note;
            16'b1000001010110000: note = 0;
            16'b1000001100010100: note = F1_note;
            16'b1000001110100110: note = 0;
            16'b1000001110111111: note = D1_note;
            16'b1000010011100011: note = 0;
            16'b1000010100010110: note = D1_note;
            16'b1000010110101000: note = 0;
            16'b1000010111000001: note = D1_note;
            16'b1000011001010011: note = 0;
            16'b1000011001101100: note = A1_note;
            16'b1000011011111110: note = 0;
            16'b1000011100010111: note = A1_note;
            16'b1000011110101001: note = 0;
            16'b1000011111000010: note = A1_note;
            16'b1000100001010100: note = 0;
            16'b1000100001101101: note = A1_note;
            16'b1000100110010001: note = 0;
            16'b1000100111000100: note = F1_note;
            16'b1000101001010110: note = 0;
            16'b1000101001101111: note = E1_note;
            16'b1000101100000001: note = 0;
            16'b1000101100011010: note = D1_note;
            16'b1000110101100011: note = 0;
            16'b1000110111000111: note = F1_note;
            16'b1000111001011001: note = 0;
            16'b1000111001110010: note = D1_note;
            16'b1000111110010110: note = 0;
            16'b1000111111001001: note = D1_note;
            16'b1001000001011011: note = 0;
            16'b1001000001110100: note = D1_note;
            16'b1001000100000110: note = 0;
            16'b1001000100011111: note = A1_note;
            16'b1001000110110001: note = 0;
            16'b1001000111001010: note = A1_note;
            16'b1001001001011100: note = 0;
            16'b1001001001110101: note = Ah1_note;
            16'b1001001100000111: note = 0;
            16'b1001001100100000: note = A2_note;
            16'b1001001101101001: note = 0;
            16'b1001001101110110: note = Ah2_note;
            16'b1001001110111111: note = 0;
            16'b1001001111001100: note = G2_note;
            16'b1001010000010101: note = 0;
            16'b1001010000100010: note = A2_note;
            16'b1001010001101011: note = 0;
            16'b1001010001111000: note = F2_note;
            16'b1001010011000001: note = 0;
            16'b1001010011001110: note = G2_note;
            16'b1001010100010111: note = 0;
            16'b1001010100100100: note = E2_note;
            16'b1001010101101101: note = 0;
            16'b1001010101111010: note = F2_note;
            16'b1001010111000011: note = 0;
            16'b1001010111010000: note = D1_note;
            16'b1001100000011001: note = 0;
            16'b1001100001111101: note = F1_note;
            16'b1001100100001111: note = 0;
            16'b1001100100101000: note = D1_note;
            16'b1001101001001100: note = 0;
            16'b1001101001111111: note = D1_note;
            16'b1001101100010001: note = 0;
            16'b1001101100101010: note = D1_note;
            16'b1001101110111100: note = 0;
            16'b1001101111010101: note = A1_note;
            16'b1001110001100111: note = 0;
            16'b1001110010000000: note = A1_note;
            16'b1001110100010010: note = 0;
            16'b1001110100101011: note = A1_note;
            16'b1001110110111101: note = 0;
            16'b1001110111010110: note = A1_note;
            16'b1001111011111010: note = 0;
            16'b1001111100101101: note = F1_note;
            16'b1001111110111111: note = 0;
            16'b1001111111011000: note = E1_note;
            16'b1010000001101010: note = 0;
            16'b1010000010000011: note = D1_note;
            16'b1010000110100111: note = 0;
            16'b1010000111011010: note = D2_note;
            16'b1010001100001110: note = 0;
            16'b1010001100110001: note = D1_note;
            16'b1010010001010101: note = 0;
            16'b1010010010001000: note = D2_note;
            16'b1010010110111100: note = 0;
            16'b1010010111011111: note = D1_note;
            16'b1010011001110001: note = 0;
            16'b1010011010001010: note = D2_note;
            16'b1010011100011100: note = 0;
            16'b1010011100110101: note = D2_note;
            16'b1010011111000111: note = 0;
            16'b1010011111100000: note = D2_note;
            16'b1010100001110010: note = 0;
            16'b1010100010001011: note = D2_note;
            16'b1010100110101111: note = 0;
            16'b1010100111100010: note = A1_note;
            16'b1010101100000110: note = 0;
            16'b1010101100111001: note = F2_note;
            16'b1010110011110000: note = 0;
            16'b1010110100111010: note = E2_note;
            16'b1010110110000011: note = 0;
            16'b1010110110010000: note = D2_note;
            16'b1010110111011001: note = 0;
            16'b1010110111100110: note = E2_note;
            16'b1010111100001010: note = 0;
            16'b1010111100111101: note = C2_note;
            16'b1011000001100001: note = 0;
            16'b1011000010010100: note = D2_note;
            16'b1011001001001011: note = 0;
            16'b1011001010010101: note = C2_note;
            16'b1011001011011110: note = 0;
            16'b1011001011101011: note = Ah1_note;
            16'b1011001100110100: note = 0;
            16'b1011001101000001: note = C2_note;
            16'b1011010001100101: note = 0;
            16'b1011010010011000: note = A1_note;
            16'b1011010110111100: note = 0;
            16'b1011010111101111: note = Ah1_note;
            16'b1011011110100110: note = 0;
            16'b1011011111110000: note = A1_note;
            16'b1011100000111001: note = 0;
            16'b1011100001000110: note = G1_note;
            16'b1011100010001111: note = 0;
            16'b1011100010011100: note = A1_note;
            16'b1011100111000000: note = 0;
            16'b1011100111110011: note = F1_note;
            16'b1011101100010111: note = 0;
            16'b1011101101001010: note = E1_note;
            16'b1011110001101110: note = 0;
            16'b1011110010100001: note = A1_note;
            16'b1011110111000101: note = 0;
            16'b1011110111111000: note = G1_note;
            16'b1011111010001010: note = 0;
            16'b1011111010100011: note = F1_note;
            16'b1011111100110101: note = 0;
            16'b1011111101001110: note = E1_note;
            16'b1011111111100000: note = 0;
            16'b1011111111111001: note = F1_note;
            16'b1100000010001011: note = 0;
            16'b1100000010100100: note = D1_note;
            16'b1100000100111101: note = 0;
            16'b1100000101010000: note = D2_note;
            16'b1100000110011001: note = 0;
            16'b1100000110100110: note = A1_note;
            16'b1100000111101111: note = 0;
            16'b1100000111111100: note = F1_note;
            16'b1100001001000101: note = 0;
            16'b1100001001010010: note = D1_note;
            16'b1100001010011011: note = 0;
            16'b1100001010101000: note = F1_note;
            16'b1100001011110001: note = 0;
            16'b1100001011111110: note = A1_note;
            16'b1100001101000111: note = 0;
            16'b1100001101010100: note = E1_note;
            16'b1100001110100000: note = 0;
            16'b1100001110101010: note = C2_note;
            16'b1100001111110011: note = 0;
            16'b1100010000000000: note = G1_note;
            16'b1100010001001001: note = 0;
            16'b1100010001010110: note = E1_note;
            16'b1100010010011111: note = 0;
            16'b1100010010101100: note = A1_note;
            16'b1100010011111000: note = 0;
            16'b1100010100000010: note = E2_note;
            16'b1100010101001011: note = 0;
            16'b1100010101011000: note = C2_note;
            16'b1100010110100001: note = 0;
            16'b1100010110101110: note = A1_note;
            16'b1100010111110111: note = 0;
            16'b1100011000000100: note = G1_note;
            16'b1100011001010000: note = 0;
            16'b1100011001011010: note = D2_note;
            16'b1100011010100011: note = 0;
            16'b1100011010110000: note = Ah1_note;
            16'b1100011011111001: note = 0;
            16'b1100011100000110: note = G1_note;
            16'b1100011101001111: note = 0;
            16'b1100011101011100: note = F2_note;
            16'b1100011110101000: note = 0;
            16'b1100011110110010: note = D3_note;
            16'b1100011111111011: note = 0;
            16'b1100100000001000: note = A2_note;
            16'b1100100001010001: note = 0;
            16'b1100100001011110: note = F2_note;
            16'b1100100010100111: note = 0;
            16'b1100100010110100: note = E2_note;
            16'b1100100101001101: note = 0;
            16'b1100100101100000: note = D2_note;
            16'b1100100111110010: note = 0;
            16'b1100101000001011: note = C2_note;
            16'b1100101010011101: note = 0;
            16'b1100101010110110: note = A1_note;
            16'b1100101101001000: note = 0;
            16'b1100101101100001: note = D2_note;
            16'b1100101110101101: note = 0;
            16'b1100101110110111: note = Ah2_note;
            16'b1100110000000000: note = 0;
            16'b1100110000001101: note = F2_note;
            16'b1100110001010110: note = 0;
            16'b1100110001100011: note = D2_note;
            16'b1100110010101100: note = 0;
            16'b1100110010111001: note = C2_note;
            16'b1100110100000101: note = 0;
            16'b1100110100001111: note = Ah2_note;
            16'b1100110101011000: note = 0;
            16'b1100110101100101: note = F2_note;
            16'b1100110110101110: note = 0;
            16'b1100110110111011: note = C2_note;
            16'b1100111000000100: note = 0;
            16'b1100111000010001: note = A1_note;
            16'b1100111001011101: note = 0;
            16'b1100111001100111: note = E2_note;
            16'b1100111010110000: note = 0;
            16'b1100111010111101: note = C2_note;
            16'b1100111100000110: note = 0;
            16'b1100111100010011: note = A1_note;
            16'b1100111101011100: note = 0;
            16'b1100111101101001: note = C2_note;
            16'b1100111110110101: note = 0;
            16'b1100111110111111: note = G2_note;
            16'b1101000000001000: note = 0;
            16'b1101000000010101: note = E2_note;
            16'b1101000001011110: note = 0;
            16'b1101000001101011: note = C2_note;
            16'b1101000010110100: note = 0;
            16'b1101000011000001: note = D2_note;
            16'b1101000111110101: note = 0;
            16'b1101001000011000: note = D3_note;
            16'b1101001001100001: note = 0;
            16'b1101001001101110: note = A2_note;
            16'b1101001010110111: note = 0;
            16'b1101001011000100: note = F2_note;
            16'b1101001100001101: note = 0;
            16'b1101001100011010: note = D2_note;
            16'b1101001101100011: note = 0;
            16'b1101001101110000: note = A2_note;
            16'b1101001110111001: note = 0;
            16'b1101001111000110: note = F2_note;
            16'b1101010000001111: note = 0;
            16'b1101010000011100: note = D2_note;
            16'b1101010001100101: note = 0;
            16'b1101010001110010: note = A1_note;
            16'b1101010010111011: note = 0;
            16'b1101010011001000: note = D2_note;
            16'b1101010100010001: note = 0;
            16'b1101010100011110: note = F2_note;
            16'b1101010101100111: note = 0;
            16'b1101010101110100: note = A2_note;
            16'b1101010110111101: note = 0;
            16'b1101010111001010: note = C3_note;
            16'b1101011000010011: note = 0;
            16'b1101011000100000: note = D2_note;
            16'b1101011101000100: note = 0;
            16'b1101011101110111: note = D2_note;
            16'b1101100010101011: note = 0;
            16'b1101100011001110: note = A1_note;
            16'b1101100101100000: note = 0;
            16'b1101100101111001: note = G1_note;
            16'b1101101000001011: note = 0;
            16'b1101101000100100: note = F1_note;
            16'b1101101101001000: note = 0;
            16'b1101101101111011: note = E1_note;
            16'b1101101111000111: note = 0;
            16'b1101101111010001: note = C2_note;
            16'b1101110000011010: note = 0;
            16'b1101110000100111: note = A1_note;
            16'b1101110001110000: note = 0;
            16'b1101110001111101: note = E1_note;
            16'b1101110011000110: note = 0;
            16'b1101110011010011: note = A1_note;
            16'b1101110100011100: note = 0;
            16'b1101110100101001: note = E1_note;
            16'b1101110101110010: note = 0;
            16'b1101110101111111: note = A1_note;
            16'b1101110111001000: note = 0;
            16'b1101110111010101: note = C2_note;
            16'b1101111000011110: note = 0;
            16'b1101111000101011: note = F1_note;
            16'b1101111101011111: note = 0;
            16'b1101111110000010: note = E1_note;
            16'b1110000000010100: note = 0;
            16'b1110000000101101: note = A2_note;
            16'b1110000001110110: note = 0;
            16'b1110000010000011: note = C3_note;
            16'b1110000011001100: note = 0;
            16'b1110000011011001: note = D2_note;
            16'b1110000111111101: note = 0;
            16'b1110001000110000: note = D3_note;
            16'b1110001101100100: note = 0;
            16'b1110001110000111: note = D2_note;
            16'b1110010010101011: note = 0;
            16'b1110010011011110: note = D3_note;
            16'b1110011000010010: note = 0;
            16'b1110011000110101: note = D2_note;
            16'b1110011011000111: note = 0;
            16'b1110011011100000: note = D3_note;
            16'b1110011101110010: note = 0;
            16'b1110011110001011: note = D3_note;
            16'b1110100000011101: note = 0;
            16'b1110100000110110: note = D3_note;
            16'b1110100011001000: note = 0;
            16'b1110100011100001: note = D3_note;
            16'b1110101100101010: note = 0;
            16'b1110101101101011: note = Dh1_note;
            16'b1110101110110111: note = 0;
            16'b1110110000010110: note = Dh1_note;
            16'b1110110001100010: note = 0;
            16'b1110110011000001: note = E1_note;
            16'b1110110100001101: note = 0;
            16'b1110110101101100: note = E1_note;
            16'b1110110110111000: note = 0;
            16'b1110111000010111: note = Dh1_note;
            16'b1110111001100011: note = 0;
            16'b1110111011000010: note = Dh1_note;
            16'b1110111100001110: note = 0;
            16'b1110111101101101: note = E1_note;
            16'b1110111110111001: note = 0;
            16'b1111000000011000: note = E1_note;
            16'b1111000001100100: note = 0;
            16'b1111000011000011: note = Dh1_note;
            16'b1111000100001111: note = 0;
            16'b1111000101101110: note = Dh1_note;
            16'b1111000110111010: note = 0;
            16'b1111001000011001: note = E1_note;
            16'b1111001001100101: note = 0;
            16'b1111001011000100: note = E1_note;
            16'b1111001100010000: note = 0;
            16'b1111001101101111: note = Dh2_note;
            16'b1111010111010111: note = 0;
            16'b1111011000011100: note = Dh1_note;
            16'b1111011001101000: note = 0;
            16'b1111011011000111: note = Dh1_note;
            16'b1111011100010011: note = 0;
            16'b1111011101110010: note = E1_note;
            16'b1111011110111110: note = 0;
            16'b1111100000011101: note = E1_note;
            16'b1111100001101001: note = 0;
            16'b1111100011001000: note = Dh1_note;
            16'b1111100100010100: note = 0;
            16'b1111100101110011: note = Dh1_note;
            16'b1111100110111111: note = 0;
            16'b1111101000011110: note = E1_note;
            16'b1111101001101010: note = 0;
            16'b1111101011001001: note = E1_note;
            16'b1111101100010101: note = 0;
            16'b1111101101110100: note = Dh1_note;
            16'b1111101111000000: note = 0;
            16'b1111110000011111: note = Dh1_note;
            16'b1111110001101011: note = 0;
            16'b1111110011001010: note = E1_note;
            16'b1111110100010110: note = 0;
            16'b1111110101110101: note = E1_note;
            16'b1111110111000001: note = 0;
            16'b1111111000100000: note = Dh2_note;
            17'b10000000010001000: note = 0;
            17'b10000000011001101: note = Dh1_note;
            17'b10000000100011001: note = 0;
            17'b10000000101111000: note = Dh1_note;
            17'b10000000111000100: note = 0;
            17'b10000001000100011: note = E1_note;
            17'b10000001001101111: note = 0;
            17'b10000001011001110: note = E1_note;
            17'b10000001100011010: note = 0;
            17'b10000001101111001: note = Dh1_note;
            17'b10000001111000101: note = 0;
            17'b10000010000100100: note = Dh1_note;
            17'b10000010001110000: note = 0;
            17'b10000010011001111: note = E1_note;
            17'b10000010100011011: note = 0;
            17'b10000010101111010: note = E1_note;
            17'b10000010111000110: note = 0;
            17'b10000011000100101: note = Dh1_note;
            17'b10000011001110001: note = 0;
            17'b10000011011010000: note = Dh1_note;
            17'b10000011100011100: note = 0;
            17'b10000011101111011: note = E1_note;
            17'b10000011111000111: note = 0;
            17'b10000100000100110: note = E1_note;
            17'b10000100001110010: note = 0;
            17'b10000100011010001: note = Dh2_note;
            17'b10000101100111001: note = 0;
            17'b10000101101111110: note = A1_note;
            17'b10000101111001010: note = 0;
            17'b10000110000101001: note = Gh1_note;
            17'b10000110001110101: note = 0;
            17'b10000110011010100: note = Fh1_note;
            17'b10000110100100000: note = 0;
            17'b10000110101111111: note = Gh1_note;
            17'b10000110111001011: note = 0;
            17'b10000111000101010: note = Fh1_note;
            17'b10000111001110110: note = 0;
            17'b10000111011010101: note = E1_note;
            17'b10000111100100001: note = 0;
            17'b10000111110000000: note = Fh1_note;
            17'b10000111111001100: note = 0;
            17'b10001000000101011: note = E1_note;
            17'b10001000001110111: note = 0;
            17'b10001000011010110: note = Dh1_note;
            17'b10001000100100010: note = 0;
            17'b10001000110000001: note = E1_note;
            17'b10001000111001101: note = 0;
            17'b10001001000101100: note = Dh1_note;
            17'b10001001001111000: note = 0;
            17'b10001001011010111: note = Ch1_note;
            17'b10001001100100011: note = 0;
            17'b10001001110000010: note = Dh1_note;
            17'b10001001111001110: note = 0;
            17'b10001010000101101: note = C1_note;
            17'b10001010001111001: note = 0;
            17'b10001010011011000: note = Ch1_note;
            17'b10001010100100100: note = 0;
            17'b10001011000101111: note = Ch1_note;
            17'b10001011011000001: note = 0;
            17'b10001011011011010: note = Ch1_note;
            17'b10001011101101100: note = 0;
            17'b10001011110000101: note = Gh2_note;
            17'b10001100000010111: note = 0;
            17'b10001100000110000: note = Ch3_note;
            17'b10001100011000010: note = 0;
            17'b10001100011011011: note = Gh3_note;
            17'b10001100101101101: note = 0;
            17'b10001100110000110: note = Ch3_note;
            17'b10001101000011000: note = 0;
            17'b10001101000110001: note = Gh2_note;
            17'b10001101011000011: note = 0;
            17'b10001101011011100: note = Ch3_note;
            17'b10001101101101110: note = 0;
            17'b10001101110000111: note = Gh3_note;
            17'b10001110000011001: note = 0;
            17'b10001110000110010: note = Ch3_note;
            17'b10001110011000100: note = 0;
            17'b10001110011011101: note = Gh2_note;
            17'b10001110101101111: note = 0;
            17'b10001110110001000: note = Ch3_note;
            17'b10001111000011010: note = 0;
            17'b10001111000110011: note = Gh3_note;
            17'b10001111011000101: note = 0;
            17'b10001111011011110: note = Ch3_note;
            17'b10001111101110000: note = 0;
            17'b10001111110001001: note = Gh2_note;
            17'b10010000000011011: note = 0;
            17'b10010000000110100: note = Ch3_note;
            17'b10010000011000110: note = 0;
            17'b10010000011011111: note = Ch1_note;
            17'b10010000101110001: note = 0;
            17'b10010000110001010: note = Ch1_note;
            17'b10010001000011100: note = 0;
            17'b10010001000110101: note = Gh2_note;
            17'b10010001011000111: note = 0;
            17'b10010001011100000: note = Ch3_note;
            17'b10010001101110010: note = 0;
            17'b10010001110001011: note = Gh3_note;
            17'b10010010000011101: note = 0;
            17'b10010010000110110: note = Ch3_note;
            17'b10010010011001000: note = 0;
            17'b10010010011100001: note = Gh2_note;
            17'b10010010101110011: note = 0;
            17'b10010010110001100: note = Ch3_note;
            17'b10010011000011110: note = 0;
            17'b10010011000110111: note = Gh3_note;
            17'b10010011011001001: note = 0;
            17'b10010011011100010: note = Ch3_note;
            17'b10010011101110100: note = 0;
            17'b10010011110001101: note = Gh2_note;
            17'b10010100000011111: note = 0;
            17'b10010100000111000: note = Ch3_note;
            17'b10010100011001010: note = 0;
            17'b10010100011100011: note = Gh3_note;
            17'b10010100101110101: note = 0;
            17'b10010100110001110: note = Ch3_note;
            17'b10010101000100000: note = 0;
            17'b10010101000111001: note = Gh2_note;
            17'b10010101011001011: note = 0;
            17'b10010101011100100: note = Ch3_note;
            17'b10010101101110110: note = 0;
            17'b10010101110001111: note = Ch1_note;
            17'b10010110000100001: note = 0;
            17'b10010110000111010: note = Ch1_note;
            17'b10010110011001100: note = 0;
            17'b10010110011100101: note = Gh2_note;
            17'b10010110101110111: note = 0;
            17'b10010110110010000: note = Ch3_note;
            17'b10010111000100010: note = 0;
            17'b10010111000111011: note = Gh3_note;
            17'b10010111011001101: note = 0;
            17'b10010111011100110: note = Ch3_note;
            17'b10010111101111000: note = 0;
            17'b10010111110010001: note = Gh2_note;
            17'b10011000000100011: note = 0;
            17'b10011000000111100: note = Ch3_note;
            17'b10011000011001110: note = 0;
            17'b10011000011100111: note = Gh3_note;
            17'b10011000101111001: note = 0;
            17'b10011000110010010: note = Ch3_note;
            17'b10011001000100100: note = 0;
            17'b10011001000111101: note = Gh2_note;
            17'b10011001011001111: note = 0;
            17'b10011001011101000: note = Ch3_note;
            17'b10011001101111010: note = 0;
            17'b10011001110010011: note = Gh3_note;
            17'b10011010000100101: note = 0;
            17'b10011010000111110: note = Ch3_note;
            17'b10011010011010000: note = 0;
            17'b10011010011101001: note = Gh2_note;
            17'b10011010101111011: note = 0;
            17'b10011010110010100: note = Ch3_note;
            17'b10011011000100110: note = 0;
            17'b10011011000111111: note = Ch1_note;
            17'b10011011011010001: note = 0;
            17'b10011011011101010: note = Ch1_note;
            17'b10011011101111100: note = 0;
            17'b10011011110010101: note = Gh2_note;
            17'b10011100000100111: note = 0;
            17'b10011100001000000: note = Ch3_note;
            17'b10011100011010010: note = 0;
            17'b10011100011101011: note = Gh3_note;
            17'b10011100101111101: note = 0;
            17'b10011100110010110: note = Ch3_note;
            17'b10011101000101000: note = 0;
            17'b10011101001000001: note = Gh2_note;
            17'b10011101011010011: note = 0;
            17'b10011101011101100: note = Ch3_note;
            17'b10011101101111110: note = 0;
            17'b10011101110010111: note = Gh3_note;
            17'b10011110000101001: note = 0;
            17'b10011110001000010: note = Ch3_note;
            17'b10011110011010100: note = 0;
            17'b10011110011101101: note = Gh2_note;
            17'b10011110101111111: note = 0;
            17'b10011110110011000: note = Ch3_note;
            17'b10011111000101010: note = 0;
            17'b10011111001000011: note = Gh3_note;
            17'b10011111011010101: note = 0;
            17'b10011111011101110: note = Ch3_note;
            17'b10011111110000000: note = 0;
            17'b10011111110011001: note = Gh2_note;
            17'b10100000000101011: note = 0;
            17'b10100000001000100: note = Ch3_note;
            17'b10100000011010110: note = 0;
            17'b10100000011101111: note = Ch1_note;
            17'b10100000110000001: note = 0;
            17'b10100000110011010: note = Ch1_note;
            17'b10100001000101100: note = 0;
            17'b10100001001000101: note = E1_note;
            17'b10100001011010111: note = 0;
            17'b10100001011110000: note = Dh1_note;
            17'b10100010000010100: note = 0;
            17'b10100010001000111: note = B_note;
            17'b10100010101101011: note = 0;
            17'b10100010110011110: note = Ch1_note;
            17'b10100101011000011: note = 0;
            17'b10100101110100011: note = Ch1_note;
            17'b10100110000110101: note = 0;
            17'b10100110001001110: note = Ch1_note;
            17'b10100110011100000: note = 0;
            17'b10100110011111001: note = E1_note;
            17'b10100110110001011: note = 0;
            17'b10100110110100100: note = Dh1_note;
            17'b10100111011001000: note = 0;
            17'b10100111011111011: note = B_note;
            17'b10101000000011111: note = 0;
            17'b10101000001010010: note = Ch1_note;
            17'b10101010101110111: note = 0;
            17'b10101011001010111: note = Ch1_note;
            17'b10101011011101001: note = 0;
            17'b10101011100000010: note = Ch1_note;
            17'b10101011110010100: note = 0;
            17'b10101011110101101: note = E1_note;
            17'b10101100000111111: note = 0;
            17'b10101100001011000: note = Dh1_note;
            17'b10101100101111100: note = 0;
            17'b10101100110101111: note = B_note;
            17'b10101101011010011: note = 0;
            17'b10101101100000110: note = Ch1_note;
            17'b10110000000101011: note = 0;
            17'b10110000010111101: note = C1_note;
            17'b10110000101001111: note = 0;
            17'b10110000101101000: note = C1_note;
            17'b10110000111111010: note = 0;
            17'b10110001000010011: note = Dh1_note;
            17'b10110001010100101: note = 0;
            17'b10110001010111110: note = Ch1_note;
            17'b10110001111100010: note = 0;
            17'b10110010000010101: note = C1_note;
            17'b10110010100111001: note = 0;
            17'b10110010101101100: note = Gh1_note;
            17'b10110011010010000: note = 0;
            17'b10110100011000101: note = Ch3_note;
            17'b10110100100001110: note = 0;
            17'b10110100100011011: note = Ch2_note;
            17'b10110100101100100: note = 0;
            17'b10110100101110001: note = B2_note;
            17'b10110100110111010: note = 0;
            17'b10110100111000111: note = B1_note;
            17'b10110101000010000: note = 0;
            17'b10110101000011101: note = A2_note;
            17'b10110101001100110: note = 0;
            17'b10110101001110011: note = A1_note;
            17'b10110101010111100: note = 0;
            17'b10110101011001001: note = Gh2_note;
            17'b10110101100010010: note = 0;
            17'b10110101100011111: note = Gh1_note;
            17'b10110101101101000: note = 0;
            17'b10110101101110101: note = Ch1_note;
            17'b10110110010101001: note = 0;
            17'b10110110011001011: note = E1_note;
            17'b10110110111100000: note = 0;
            17'b10110111000100010: note = E1_note;
            17'b10110111010110100: note = 0;
            17'b10110111011001101: note = Ch1_note;
            17'b10110111111110001: note = 0;
            17'b10111000000100100: note = Ch1_note;
            17'b10111000010110110: note = 0;
            17'b10111000011001111: note = Ch1_note;
            17'b10111000101100001: note = 0;
            17'b10111000101111010: note = Gh1_note;
            17'b10111001000001100: note = 0;
            17'b10111001000100101: note = Gh1_note;
            17'b10111001010110111: note = 0;
            17'b10111001011010000: note = Gh1_note;
            17'b10111001101100010: note = 0;
            17'b10111001101111011: note = Gh1_note;
            17'b10111010010011111: note = 0;
            17'b10111010011010010: note = E1_note;
            17'b10111010101100100: note = 0;
            17'b10111010101111101: note = Dh1_note;
            17'b10111011000001111: note = 0;
            17'b10111011000101000: note = Ch1_note;
            17'b10111100001110001: note = 0;
            17'b10111100011010101: note = E1_note;
            17'b10111100101100111: note = 0;
            17'b10111100110000000: note = Ch1_note;
            17'b10111101010100100: note = 0;
            17'b10111101011010111: note = Ch1_note;
            17'b10111101101101001: note = 0;
            17'b10111101110000010: note = Ch1_note;
            17'b10111110000010100: note = 0;
            17'b10111110000101101: note = Gh1_note;
            17'b10111110010111111: note = 0;
            17'b10111110011011000: note = Gh1_note;
            17'b10111110101101010: note = 0;
            17'b10111110110000011: note = Gh1_note;
            17'b10111111000010101: note = 0;
            17'b10111111000101110: note = Ch2_note;
            17'b10111111011000000: note = 0;
            17'b10111111011011001: note = B1_note;
            17'b10111111101101011: note = 0;
            17'b10111111110000100: note = A1_note;
            17'b11000000000010110: note = 0;
            17'b11000000000101111: note = Gh1_note;
            17'b11000000011000001: note = 0;
            17'b11000000011011010: note = Ch1_note;
            17'b11000001000001110: note = 0;
            17'b11000001000110000: note = E1_note;
            17'b11000001101000101: note = 0;
            17'b11000001110000111: note = E1_note;
            17'b11000010000011001: note = 0;
            17'b11000010000110010: note = Ch1_note;
            17'b11000010101010110: note = 0;
            17'b11000010110001001: note = Ch1_note;
            17'b11000011000011011: note = 0;
            17'b11000011000110100: note = Ch1_note;
            17'b11000011011000110: note = 0;
            17'b11000011011011111: note = Gh1_note;
            17'b11000011101110001: note = 0;
            17'b11000011110001010: note = Gh1_note;
            17'b11000100000011100: note = 0;
            17'b11000100000110101: note = Gh1_note;
            17'b11000100011000111: note = 0;
            17'b11000100011100000: note = Gh1_note;
            17'b11000101000000100: note = 0;
            17'b11000101000110111: note = E1_note;
            17'b11000101011001001: note = 0;
            17'b11000101011100010: note = Dh1_note;
            17'b11000101101110100: note = 0;
            17'b11000101110001101: note = Ch1_note;
            17'b11000110010110001: note = 0;
            17'b11000110011100100: note = Ch2_note;
            17'b11000111000011000: note = 0;
            17'b11000111000111011: note = Ch1_note;
            17'b11000111101011111: note = 0;
            17'b11000111110010010: note = Ch2_note;
            17'b11001000011000110: note = 0;
            17'b11001000011101001: note = Ch1_note;
            17'b11001000101111011: note = 0;
            17'b11001000110010100: note = Ch2_note;
            17'b11001001000100110: note = 0;
            17'b11001001000111111: note = Ch2_note;
            17'b11001001011010001: note = 0;
            17'b11001001011101010: note = Ch2_note;
            17'b11001001101111100: note = 0;
            17'b11001001110010101: note = Ch2_note;
            17'b11001010000100111: note = 0;
            17'b11001010001000000: note = B1_note;
            17'b11001010011010010: note = 0;
            17'b11001010011101011: note = A1_note;
            17'b11001010101111101: note = 0;
            17'b11001010110010110: note = Ch2_note;
            17'b11001010111011111: note = 0;
            17'b11001010111101100: note = Dh2_note;
            17'b11001011000110101: note = 0;
            17'b11001011001000010: note = E2_note;
            17'b11001011011010100: note = 0;
            17'b11001011011101101: note = Dh2_note;
            17'b11001011101111111: note = 0;
            17'b11001011110011000: note = Fh2_note;
            17'b11001100000101010: note = 0;
            17'b11001100001000011: note = E2_note;
            17'b11001100011010101: note = 0;
            17'b11001100011101110: note = Gh2_note;
            17'b11001100110000000: note = 0;
            17'b11001100110011001: note = Fh2_note;
            17'b11001101000101011: note = 0;
            17'b11001101001000100: note = A2_note;
            17'b11001101011010110: note = 0;
            17'b11001101011101111: note = Gh2_note;
            17'b11001101110000001: note = 0;
            17'b11001101110011010: note = Fh2_note;
            17'b11001110000101100: note = 0;
            17'b11001110001000101: note = Gh2_note;
            17'b11001110011010111: note = 0;
            17'b11001110011110000: note = E2_note;
            17'b11001110110000010: note = 0;
            17'b11001110110011011: note = Dh2_note;
            17'b11001111000101101: note = 0;
            17'b11001111001000110: note = E2_note;
            17'b11001111011011000: note = 0;
            17'b11001111011110001: note = Gh2_note;
            17'b11001111110000011: note = 0;
            17'b11001111110011100: note = Dh2_note;
            17'b11010000000101110: note = 0;
            17'b11010000001000111: note = Gh2_note;
            17'b11010000011011001: note = 0;
            17'b11010000011110010: note = Ch2_note;
            17'b11010000110000100: note = 0;
            17'b11010000110011101: note = Gh1_note;
            17'b11010001000101111: note = 0;
            17'b11010001001001000: note = Ch2_note;
            17'b11010001011011010: note = 0;
            17'b11010001011110011: note = Dh2_note;
            17'b11010001110000101: note = 0;
            17'b11010001110011110: note = E2_note;
            17'b11010010000110000: note = 0;
            17'b11010010001001001: note = Gh1_note;
            17'b11010010011011011: note = 0;
            17'b11010010011110100: note = Dh2_note;
            17'b11010010110000110: note = 0;
            17'b11010010110011111: note = Gh1_note;
            17'b11010011000110001: note = 0;
            17'b11010011001001010: note = Ch2_note;
            17'b11010011011011100: note = 0;
            17'b11010011011110101: note = Gh1_note;
            17'b11010011110000111: note = 0;
            17'b11010011110100000: note = Ch2_note;
            17'b11010100000110010: note = 0;
            17'b11010100001001011: note = Gh1_note;
            17'b11010100011011101: note = 0;
            17'b11010100011110110: note = Ch2_note;
            17'b11010100110001000: note = 0;
            17'b11010100110100001: note = B1_note;
            17'b11010101000110011: note = 0;
            17'b11010101001001100: note = Gh2_note;
            17'b11010101101110000: note = 0;
            17'b11010101110100011: note = E3_note;
            17'b11010110011000111: note = 0;
            17'b11010110011111010: note = Fh3_note;
            17'b11010110110001100: note = 0;
            17'b11010110110100101: note = Dh3_note;
            17'b11010111011001001: note = 0;
            17'b11010111011111100: note = E3_note;
            17'b11011000000100000: note = 0;
            17'b11011000001010011: note = Ch3_note;
            17'b11011000101110111: note = 0;
            17'b11011000110101010: note = Dh3_note;
            17'b11011001011001110: note = 0;
            17'b11011001100000001: note = A2_note;
            17'b11011010000100101: note = 0;
            17'b11011010001011000: note = Gh2_note;
            17'b11011010101111100: note = 0;
            17'b11011010110101111: note = Gh2_note;
            17'b11011011001000001: note = 0;
            17'b11011011001011010: note = E3_note;
            17'b11011011101111110: note = 0;
            17'b11011011110110001: note = Fh3_note;
            17'b11011100001000011: note = 0;
            17'b11011100001011100: note = Dh3_note;
            17'b11011100110000000: note = 0;
            17'b11011100110110011: note = E3_note;
            17'b11011101011010111: note = 0;
            17'b11011101100001010: note = Ch3_note;
            17'b11011110000101110: note = 0;
            17'b11011110001100001: note = B3_note;
            17'b11011110110000101: note = 0;
            17'b11011110110111000: note = Ch4_note;
            17'b11011111101101111: note = 0;
            17'b11011111110111001: note = Gh2_note;
            17'b11100000011011101: note = 0;
            17'b11100000100010000: note = E3_note;
            17'b11100001000110100: note = 0;
            17'b11100001001100111: note = Fh3_note;
            17'b11100001011111001: note = 0;
            17'b11100001100010010: note = Dh3_note;
            17'b11100010000110110: note = 0;
            17'b11100010001101001: note = E3_note;
            17'b11100010110001101: note = 0;
            17'b11100010111000000: note = Ch3_note;
            17'b11100011011100100: note = 0;
            17'b11100011100010111: note = Dh3_note;
            17'b11100100000111011: note = 0;
            17'b11100100001101110: note = A2_note;
            17'b11100100110010010: note = 0;
            17'b11100100111000101: note = Gh2_note;
            17'b11100101101111100: note = 0;
            17'b11100101111000110: note = E2_note;
            17'b11100110011101010: note = 0;
            17'b11100110100011101: note = Gh2_note;
            17'b11100110110101111: note = 0;
            17'b11100110111001000: note = Dh2_note;
            17'b11100111011101100: note = 0;
            17'b11100111100011111: note = Gh2_note;
            17'b11101000001000011: note = 0;
            17'b11101000001110110: note = E1_note;
            17'b11101000100001000: note = 0;
            17'b11101001111000101: note = D3_note;
            17'b11101010000001110: note = 0;
            17'b11101010000011011: note = D2_note;
            17'b11101010001100100: note = 0;
            17'b11101010001110001: note = C3_note;
            17'b11101010010111010: note = 0;
            17'b11101010011000111: note = C2_note;
            17'b11101010100010000: note = 0;
            17'b11101010100011101: note = Ah2_note;
            17'b11101010101100110: note = 0;
            17'b11101010101110011: note = Ah1_note;
            17'b11101010110111100: note = 0;
            17'b11101010111001001: note = A2_note;
            17'b11101011000010010: note = 0;
            17'b11101011000011111: note = A1_note;
            17'b11101011001101000: note = 0;
            17'b11101011001110101: note = D1_note;
            17'b11101100010111110: note = 0;
            17'b11101100100100010: note = F1_note;
            17'b11101100110110100: note = 0;
            17'b11101100111001101: note = D1_note;
            17'b11101101011110001: note = 0;
            17'b11101101100100100: note = D1_note;
            17'b11101101110110110: note = 0;
            17'b11101101111001111: note = D1_note;
            17'b11101110001100001: note = 0;
            17'b11101110001111010: note = A1_note;
            17'b11101110100001100: note = 0;
            17'b11101110100100101: note = A1_note;
            17'b11101110110110111: note = 0;
            17'b11101110111010000: note = A1_note;
            17'b11101111001100010: note = 0;
            17'b11101111001111011: note = A1_note;
            17'b11101111110011111: note = 0;
            17'b11101111111010010: note = F1_note;
            17'b11110000001100100: note = 0;
            17'b11110000001111101: note = E1_note;
            17'b11110000100001111: note = 0;
            17'b11110000100101000: note = D1_note;
            17'b11110001101110001: note = 0;
            17'b11110001111010101: note = F1_note;
            17'b11110010001100111: note = 0;
            17'b11110010010000000: note = D1_note;
            17'b11110010110100100: note = 0;
            17'b11110010111010111: note = D1_note;
            17'b11110011001101001: note = 0;
            17'b11110011010000010: note = D1_note;
            17'b11110011100010100: note = 0;
            17'b11110011100101101: note = A1_note;
            17'b11110011110111111: note = 0;
            17'b11110011111011000: note = A1_note;
            17'b11110100001101010: note = 0;
            17'b11110100010000011: note = Ah1_note;
            17'b11110100100010101: note = 0;
            17'b11110100100101110: note = A2_note;
            17'b11110100101110111: note = 0;
            17'b11110100110000100: note = Ah2_note;
            17'b11110100111001101: note = 0;
            17'b11110100111011010: note = G2_note;
            17'b11110101000100011: note = 0;
            17'b11110101000110000: note = A2_note;
            17'b11110101001111001: note = 0;
            17'b11110101010000110: note = F2_note;
            17'b11110101011001111: note = 0;
            17'b11110101011011100: note = G2_note;
            17'b11110101100100101: note = 0;
            17'b11110101100110010: note = E2_note;
            17'b11110101101111011: note = 0;
            17'b11110101110001000: note = F2_note;
            17'b11110101111010001: note = 0;
            17'b11110101111011110: note = D1_note;
            17'b11110111000100111: note = 0;
            17'b11110111010001011: note = F1_note;
            17'b11110111100011101: note = 0;
            17'b11110111100110110: note = D1_note;
            17'b11111000001011010: note = 0;
            17'b11111000010001101: note = D1_note;
            17'b11111000100011111: note = 0;
            17'b11111000100111000: note = D1_note;
            17'b11111000111001010: note = 0;
            17'b11111000111100011: note = A1_note;
            17'b11111001001110101: note = 0;
            17'b11111001010001110: note = A1_note;
            17'b11111001100100000: note = 0;
            17'b11111001100111001: note = A1_note;
            17'b11111001111001011: note = 0;
            17'b11111001111100100: note = A1_note;
            17'b11111010100001000: note = 0;
            17'b11111010100111011: note = F1_note;
            17'b11111010111001101: note = 0;
            17'b11111010111100110: note = E1_note;
            17'b11111011001111000: note = 0;
            17'b11111011010010001: note = D1_note;
            17'b11111011110110101: note = 0;
            17'b11111011111101000: note = D2_note;
            17'b11111100100011100: note = 0;
            17'b11111100100111111: note = D1_note;
            17'b11111101001100011: note = 0;
            17'b11111101010010110: note = D2_note;
            17'b11111101111001010: note = 0;
            17'b11111101111101101: note = D1_note;
            17'b11111110001111111: note = 0;
            17'b11111110010011000: note = D2_note;
            17'b11111110100101010: note = 0;
            17'b11111110101000011: note = D2_note;
            17'b11111110111010101: note = 0;
            17'b11111110111101110: note = D2_note;
            17'b11111111010000000: note = 0;
            17'b11111111010011001: note = D2_note;
            17'b11111111110111101: note = 0;
            17'b11111111111110000: note = A1_note;
            18'b100000000100010100: note = 0;
            18'b100000000101000111: note = D1_note;
            18'b100000000111011001: note = 0;
            18'b100000000111110010: note = A1_note;
            18'b100000001100010110: note = 0;
            18'b100000001101001001: note = Ah1_note;
            18'b100000010001101101: note = 0;
            18'b100000010010100000: note = G1_note;
            18'b100000010111000100: note = 0;
            18'b100000010111110111: note = A1_note;
            18'b100000011010001001: note = 0;
            18'b100000011010100010: note = D1_note;
            18'b100000011100110100: note = 0;
            18'b100000011101001101: note = A1_note;
            18'b100000100001110001: note = 0;
            18'b100000100010100100: note = Ah1_note;
            18'b100000100111001000: note = 0;
            18'b100000100111111011: note = G1_note;
            18'b100000101100011111: note = 0;
            18'b100000101101010010: note = A1_note;
            18'b100000101111100100: note = 0;
            18'b100000101111111101: note = D1_note;
            18'b100000110010001111: note = 0;
            18'b100000110010101000: note = A1_note;
            18'b100000110111001100: note = 0;
            18'b100000110111111111: note = Ah1_note;
            18'b100000111100100011: note = 0;
            18'b100000111101010110: note = G1_note;
            18'b100001000001111010: note = 0;
            18'b100001000010101101: note = A1_note;
            18'b100001000111010001: note = 0;
            18'b100001001000000100: note = F1_note;
            18'b100001001100101000: note = 0;
            18'b100001001101011011: note = G1_note;
            18'b100001010001111111: note = 0;
            18'b100001010010110010: note = E1_note;
            18'b100001010111010110: note = 0;
            18'b100001011000001001: note = F1_note;
            18'b100001011010011011: note = 0;
            18'b100001011010110100: note = D1_note;
            18'b100001011101001101: note = 0;
            18'b100001011101100000: note = D2_note;
            18'b100001011110101001: note = 0;
            18'b100001011110110110: note = A1_note;
            18'b100001011111111111: note = 0;
            18'b100001100000001100: note = F1_note;
            18'b100001100001010101: note = 0;
            18'b100001100001100010: note = D1_note;
            18'b100001100010101011: note = 0;
            18'b100001100010111000: note = F1_note;
            18'b100001100100000001: note = 0;
            18'b100001100100001110: note = A1_note;
            18'b100001100101010111: note = 0;
            18'b100001100101100100: note = E1_note;
            18'b100001100110110000: note = 0;
            18'b100001100110111010: note = C2_note;
            18'b100001101000000011: note = 0;
            18'b100001101000010000: note = G1_note;
            18'b100001101001011001: note = 0;
            18'b100001101001100110: note = E1_note;
            18'b100001101010101111: note = 0;
            18'b100001101010111100: note = A1_note;
            18'b100001101100001000: note = 0;
            18'b100001101100010010: note = E2_note;
            18'b100001101101011011: note = 0;
            18'b100001101101101000: note = C2_note;
            18'b100001101110110001: note = 0;
            18'b100001101110111110: note = A1_note;
            18'b100001110000000111: note = 0;
            18'b100001110000010100: note = G1_note;
            18'b100001110001100000: note = 0;
            18'b100001110001101010: note = D2_note;
            18'b100001110010110011: note = 0;
            18'b100001110011000000: note = Ah1_note;
            18'b100001110100001001: note = 0;
            18'b100001110100010110: note = G1_note;
            18'b100001110101011111: note = 0;
            18'b100001110101101100: note = F2_note;
            18'b100001110110111000: note = 0;
            18'b100001110111000010: note = D3_note;
            18'b100001111000001011: note = 0;
            18'b100001111000011000: note = A2_note;
            18'b100001111001100001: note = 0;
            18'b100001111001101110: note = F2_note;
            18'b100001111010110111: note = 0;
            18'b100001111011000100: note = E2_note;
            18'b100001111101011101: note = 0;
            18'b100001111101110000: note = D2_note;
            18'b100010000000000010: note = 0;
            18'b100010000000011011: note = C2_note;
            18'b100010000010101101: note = 0;
            18'b100010000011000110: note = A1_note;
            18'b100010000101011000: note = 0;
            18'b100010000101110001: note = D2_note;
            18'b100010000110111101: note = 0;
            18'b100010000111000111: note = Ah2_note;
            18'b100010001000010000: note = 0;
            18'b100010001000011101: note = F2_note;
            18'b100010001001100110: note = 0;
            18'b100010001001110011: note = D2_note;
            18'b100010001010111100: note = 0;
            18'b100010001011001001: note = C2_note;
            18'b100010001100010101: note = 0;
            18'b100010001100011111: note = Ah2_note;
            18'b100010001101101000: note = 0;
            18'b100010001101110101: note = F2_note;
            18'b100010001110111110: note = 0;
            18'b100010001111001011: note = C2_note;
            18'b100010010000010100: note = 0;
            18'b100010010000100001: note = A1_note;
            18'b100010010001101101: note = 0;
            18'b100010010001110111: note = E2_note;
            18'b100010010011000000: note = 0;
            18'b100010010011001101: note = C2_note;
            18'b100010010100010110: note = 0;
            18'b100010010100100011: note = A1_note;
            18'b100010010101101100: note = 0;
            18'b100010010101111001: note = C2_note;
            18'b100010010111000101: note = 0;
            18'b100010010111001111: note = G2_note;
            18'b100010011000011000: note = 0;
            18'b100010011000100101: note = E2_note;
            18'b100010011001101110: note = 0;
            18'b100010011001111011: note = C2_note;
            18'b100010011011000100: note = 0;
            18'b100010011011010001: note = D2_note;
            18'b100010100000000101: note = 0;
            18'b100010100000101000: note = D3_note;
            18'b100010100001110001: note = 0;
            18'b100010100001111110: note = A2_note;
            18'b100010100011000111: note = 0;
            18'b100010100011010100: note = F2_note;
            18'b100010100100011101: note = 0;
            18'b100010100100101010: note = D2_note;
            18'b100010100101110011: note = 0;
            18'b100010100110000000: note = A2_note;
            18'b100010100111001001: note = 0;
            18'b100010100111010110: note = F2_note;
            18'b100010101000011111: note = 0;
            18'b100010101000101100: note = D2_note;
            18'b100010101001110101: note = 0;
            18'b100010101010000010: note = A1_note;
            18'b100010101011001011: note = 0;
            18'b100010101011011000: note = D2_note;
            18'b100010101100100001: note = 0;
            18'b100010101100101110: note = F2_note;
            18'b100010101101110111: note = 0;
            18'b100010101110000100: note = A2_note;
            18'b100010101111001101: note = 0;
            18'b100010101111011010: note = C3_note;
            18'b100010110000100011: note = 0;
            18'b100010110000110000: note = D2_note;
            18'b100010110101010100: note = 0;
            18'b100010110110000111: note = D2_note;
            18'b100010111010111011: note = 0;
            18'b100010111011011110: note = A1_note;
            18'b100010111101110000: note = 0;
            18'b100010111110001001: note = G1_note;
            18'b100011000000011011: note = 0;
            18'b100011000000110100: note = F1_note;
            18'b100011000101011000: note = 0;
            18'b100011000110001011: note = E1_note;
            18'b100011000111010111: note = 0;
            18'b100011000111100001: note = C2_note;
            18'b100011001000101010: note = 0;
            18'b100011001000110111: note = A1_note;
            18'b100011001010000000: note = 0;
            18'b100011001010001101: note = E1_note;
            18'b100011001011010110: note = 0;
            18'b100011001011100011: note = A1_note;
            18'b100011001100101100: note = 0;
            18'b100011001100111001: note = E1_note;
            18'b100011001110000010: note = 0;
            18'b100011001110001111: note = A1_note;
            18'b100011001111011000: note = 0;
            18'b100011001111100101: note = C2_note;
            18'b100011010000101110: note = 0;
            18'b100011010000111011: note = F1_note;
            18'b100011010101101111: note = 0;
            18'b100011010110010010: note = E1_note;
            18'b100011011000100100: note = 0;
            18'b100011011000111101: note = A2_note;
            18'b100011011010000110: note = 0;
            18'b100011011010010011: note = C3_note;
            18'b100011011011011100: note = 0;
            18'b100011011011101001: note = D2_note;
            18'b100011100000001101: note = 0;
            18'b100011100001000000: note = D3_note;
            18'b100011100101110100: note = 0;
            18'b100011100110010111: note = D2_note;
            18'b100011101010111011: note = 0;
            18'b100011101011101110: note = D3_note;
            18'b100011110000100010: note = 0;
            18'b100011110001000101: note = D2_note;
            18'b100011110011010111: note = 0;
            18'b100011110011110000: note = D3_note;
            18'b100011110110000010: note = 0;
            18'b100011110110011011: note = D3_note;
            18'b100011111000101101: note = 0;
            18'b100011111001000110: note = D3_note;
            18'b100011111011011000: note = 0;
            18'b100011111011110001: note = D3_note;
            18'b100100000100111010: note = 0;
            18'b100100000101111011: note = Dh1_note;
            18'b100100000111000111: note = 0;
            18'b100100001000100110: note = Dh1_note;
            18'b100100001001110010: note = 0;
            18'b100100001011010001: note = E1_note;
            18'b100100001100011101: note = 0;
            18'b100100001101111100: note = E1_note;
            18'b100100001111001000: note = 0;
            18'b100100010000100111: note = Dh1_note;
            18'b100100010001110011: note = 0;
            18'b100100010011010010: note = Dh1_note;
            18'b100100010100011110: note = 0;
            18'b100100010101111101: note = E1_note;
            18'b100100010111001001: note = 0;
            18'b100100011000101000: note = E1_note;
            18'b100100011001110100: note = 0;
            18'b100100011011010011: note = Dh1_note;
            18'b100100011100011111: note = 0;
            18'b100100011101111110: note = Dh1_note;
            18'b100100011111001010: note = 0;
            18'b100100100000101001: note = E1_note;
            18'b100100100001110101: note = 0;
            18'b100100100011010100: note = E1_note;
            18'b100100100100100000: note = 0;
            18'b100100100101111111: note = Dh2_note;
            18'b100100101111100111: note = 0;
            18'b100100110000101100: note = Dh1_note;
            18'b100100110001111000: note = 0;
            18'b100100110011010111: note = Dh1_note;
            18'b100100110100100011: note = 0;
            18'b100100110110000010: note = E1_note;
            18'b100100110111001110: note = 0;
            18'b100100111000101101: note = E1_note;
            18'b100100111001111001: note = 0;
            18'b100100111011011000: note = Dh1_note;
            18'b100100111100100100: note = 0;
        endcase    
    end  
    //rockstar
    else if (sw_state == 4'b0100) begin
        case (counter_sec) 
            2'b11: note = Ah_note;
            8'b10001110: note = 0;
            8'b10011101: note = Ah_note;
            9'b100101011: note = 0;
            9'b100111010: note = Ah_note;
            9'b111001000: note = 0;
            9'b111010111: note = Ah_note;
            10'b1001100101: note = 0;
            10'b1001110100: note = Ah_note;
            10'b1100000010: note = 0;
            10'b1100010001: note = Ah_note;
            10'b1110011111: note = 0;
            10'b1110101110: note = Ah_note;
            11'b10000111100: note = 0;
            11'b10001001011: note = Ah_note;
            11'b10011011001: note = 0;
            11'b10011101000: note = A_note;
            11'b10101110110: note = 0;
            11'b10110000101: note = A_note;
            11'b11000010011: note = 0;
            11'b11000100010: note = A_note;
            11'b11010110000: note = 0;
            11'b11010111111: note = A_note;
            11'b11101001101: note = 0;
            11'b11101011100: note = A_note;
            12'b100001110111: note = 0;
            12'b100010010110: note = Ah_note;
            12'b100100100100: note = 0;
            12'b100100110011: note = A_note;
            12'b100111000001: note = 0;
            12'b100111010000: note = G_note;
            12'b111000111100: note = 0;
            13'b1001110100100: note = Ah_note;
            13'b1010000110010: note = 0;
            13'b1010001000001: note = Ah_note;
            13'b1010011001111: note = 0;
            13'b1010011011110: note = Ah_note;
            13'b1010101101100: note = 0;
            13'b1010101111011: note = Ah_note;
            13'b1011000001001: note = 0;
            13'b1011000011000: note = Ah_note;
            13'b1011010100110: note = 0;
            13'b1011010110101: note = Ah_note;
            13'b1011101000011: note = 0;
            13'b1011101010010: note = Ah_note;
            13'b1011111100000: note = 0;
            13'b1011111101111: note = Ah_note;
            13'b1100001111101: note = 0;
            13'b1100010001100: note = A_note;
            13'b1100100011010: note = 0;
            13'b1100100101001: note = A_note;
            13'b1100110110111: note = 0;
            13'b1100111000110: note = A_note;
            13'b1101001010100: note = 0;
            13'b1101001100011: note = A_note;
            13'b1101011110001: note = 0;
            13'b1101100000000: note = A_note;
            13'b1110000011011: note = 0;
            13'b1110000111010: note = Ah_note;
            13'b1110011001000: note = 0;
            13'b1110011010111: note = A_note;
            13'b1110101100101: note = 0;
            13'b1110101110100: note = G_note;
            14'b10000111100000: note = 0;
            14'b10011101001000: note = Ah_note;
            14'b10011111010110: note = 0;
            14'b10011111100101: note = Ah_note;
            14'b10100001110011: note = 0;
            14'b10100010000010: note = Ah_note;
            14'b10100100010000: note = 0;
            14'b10100100011111: note = Ah_note;
            14'b10100110101101: note = 0;
            14'b10100110111100: note = Ah_note;
            14'b10101001001010: note = 0;
            14'b10101001011001: note = Ah_note;
            14'b10101011100111: note = 0;
            14'b10101011110110: note = Ah_note;
            14'b10101110000100: note = 0;
            14'b10101110010011: note = Ah_note;
            14'b10110000100001: note = 0;
            14'b10110000110000: note = A_note;
            14'b10110010111110: note = 0;
            14'b10110011001101: note = A_note;
            14'b10110101011011: note = 0;
            14'b10110101101010: note = A_note;
            14'b10110111111000: note = 0;
            14'b10111000000111: note = A_note;
            14'b10111010010101: note = 0;
            14'b10111010100100: note = A_note;
            14'b10111110111111: note = 0;
            14'b10111111011110: note = Ah_note;
            14'b11000001101100: note = 0;
            14'b11000001111011: note = A_note;
            14'b11000100001001: note = 0;
            14'b11000100011000: note = G_note;
            14'b11010110000100: note = 0;
            14'b11101011101100: note = Ah_note;
            14'b11101101111010: note = 0;
            14'b11101110001001: note = Ah_note;
            14'b11110000010111: note = 0;
            14'b11110000100110: note = Ah_note;
            14'b11110010110100: note = 0;
            14'b11110011000011: note = Ah_note;
            14'b11110101010001: note = 0;
            14'b11110101100000: note = Ah_note;
            14'b11110111101110: note = 0;
            14'b11110111111101: note = Ah_note;
            14'b11111010001011: note = 0;
            14'b11111010011010: note = Ah_note;
            14'b11111100101000: note = 0;
            14'b11111100110111: note = Ah_note;
            14'b11111111000101: note = 0;
            14'b11111111010100: note = A_note;
            15'b100000001100010: note = 0;
            15'b100000001110001: note = A_note;
            15'b100000011111111: note = 0;
            15'b100000100001110: note = A_note;
            15'b100000110011100: note = 0;
            15'b100000110101011: note = A_note;
            15'b100001000111001: note = 0;
            15'b100001001001000: note = A_note;
            15'b100001101100011: note = 0;
            15'b100001110000010: note = Ah_note;
            15'b100010000010000: note = 0;
            15'b100010000011111: note = A_note;
            15'b100010010101101: note = 0;
            15'b100010010111100: note = G_note;
            15'b100100100101000: note = 0;
            15'b100111010010000: note = Ah_note;
            15'b100111100011110: note = 0;
            15'b100111100101101: note = Ah_note;
            15'b100111110111011: note = 0;
            15'b100111111001010: note = Ah_note;
            15'b101000001011000: note = 0;
            15'b101000001100111: note = Ah_note;
            15'b101000011110101: note = 0;
            15'b101000100000100: note = Ah_note;
            15'b101000110010010: note = 0;
            15'b101000110100001: note = Ah_note;
            15'b101001000101111: note = 0;
            15'b101001000111110: note = Ah_note;
            15'b101001011001100: note = 0;
            15'b101001011011011: note = Ah_note;
            15'b101001101101001: note = 0;
            15'b101001101111000: note = A_note;
            15'b101010000000110: note = 0;
            15'b101010000010101: note = A_note;
            15'b101010010100011: note = 0;
            15'b101010010110010: note = A_note;
            15'b101010101000000: note = 0;
            15'b101010101001111: note = A_note;
            15'b101010111011101: note = 0;
            15'b101010111101100: note = A_note;
            15'b101011100000111: note = 0;
            15'b101011100100110: note = Ah_note;
            15'b101011110110100: note = 0;
            15'b101011111000011: note = A_note;
            15'b101100001010001: note = 0;
            15'b101100001100000: note = G_note;
            15'b101110011001100: note = 0;
            15'b110001000110100: note = Ah_note;
            15'b110001011000010: note = 0;
            15'b110001011010001: note = Ah_note;
            15'b110001101011111: note = 0;
            15'b110001101101110: note = Ah_note;
            15'b110001111111100: note = 0;
            15'b110010000001011: note = Ah_note;
            15'b110010010011001: note = 0;
            15'b110010010101000: note = Ah_note;
            15'b110010100110110: note = 0;
            15'b110010101000101: note = Ah_note;
            15'b110010111010011: note = 0;
            15'b110010111100010: note = Ah_note;
            15'b110011001110000: note = 0;
            15'b110011001111111: note = Ah_note;
            15'b110011100001101: note = 0;
            15'b110011100011100: note = A_note;
            15'b110011110101010: note = 0;
            15'b110011110111001: note = A_note;
            15'b110100001000111: note = 0;
            15'b110100001010110: note = A_note;
            15'b110100011100100: note = 0;
            15'b110100011110011: note = A_note;
            15'b110100110000001: note = 0;
            15'b110100110010000: note = A_note;
            15'b110101010101011: note = 0;
            15'b110101011001010: note = Ah_note;
            15'b110101101011000: note = 0;
            15'b110101101100111: note = A_note;
            15'b110101111110101: note = 0;
            15'b110110000000100: note = G_note;
            15'b111000001110000: note = 0;
            15'b111010111011000: note = Ah_note;
            15'b111011001100110: note = 0;
            15'b111011001110101: note = Ah_note;
            15'b111011100000011: note = 0;
            15'b111011100010010: note = Ah_note;
            15'b111011110100000: note = 0;
            15'b111011110101111: note = Ah_note;
            15'b111100000111101: note = 0;
            15'b111100001001100: note = Ah_note;
            15'b111100011011010: note = 0;
            15'b111100011101001: note = Ah_note;
            15'b111100101110111: note = 0;
            15'b111100110000110: note = Ah_note;
            15'b111101000010100: note = 0;
            15'b111101000100011: note = Ah_note;
            15'b111101010110001: note = 0;
            15'b111101011000000: note = A_note;
            15'b111101101001110: note = 0;
            15'b111101101011101: note = A_note;
            15'b111101111101011: note = 0;
            15'b111101111111010: note = A_note;
            15'b111110010001000: note = 0;
            15'b111110010010111: note = A_note;
            15'b111110100100101: note = 0;
            15'b111110100110100: note = A_note;
            15'b111111001001111: note = 0;
            15'b111111001101110: note = Ah_note;
            15'b111111011111100: note = 0;
            15'b111111100001011: note = A_note;
            15'b111111110011001: note = 0;
            15'b111111110101000: note = G_note;
            16'b1000010000010100: note = 0;
            16'b1000100101111100: note = Ah_note;
            16'b1000101000001010: note = 0;
            16'b1000101000011001: note = Ah_note;
            16'b1000101010100111: note = 0;
            16'b1000101010110110: note = Ah_note;
            16'b1000101101000100: note = 0;
            16'b1000101101010011: note = Ah_note;
            16'b1000101111100001: note = 0;
            16'b1000101111110000: note = Ah_note;
            16'b1000110001111110: note = 0;
            16'b1000110010001101: note = Ah_note;
            16'b1000110100011011: note = 0;
            16'b1000110100101010: note = Ah_note;
            16'b1000110110111000: note = 0;
            16'b1000110111000111: note = Ah_note;
            16'b1000111001010101: note = 0;
            16'b1000111001100100: note = A_note;
            16'b1000111011110010: note = 0;
            16'b1000111100000001: note = A_note;
            16'b1000111110001111: note = 0;
            16'b1000111110011110: note = A_note;
            16'b1001000000101100: note = 0;
            16'b1001000000111011: note = A_note;
            16'b1001000011001001: note = 0;
            16'b1001000011011000: note = A_note;
            16'b1001000111110011: note = 0;
            16'b1001001000010010: note = Ah_note;
            16'b1001001010100000: note = 0;
            16'b1001001010101111: note = A_note;
            16'b1001001100111101: note = 0;
            16'b1001010010000110: note = D1_note;
            16'b1001010100010100: note = 0;
            16'b1001010100100011: note = D1_note;
            16'b1001010110110001: note = 0;
            16'b1001010111000000: note = D1_note;
            16'b1001011001001110: note = 0;
            16'b1001011001011101: note = D1_note;
            16'b1001011011101011: note = 0;
            16'b1001011011111010: note = D1_note;
            16'b1001011110001000: note = 0;
            16'b1001011110010111: note = D1_note;
            16'b1001100000100101: note = 0;
            16'b1001100000110100: note = D1_note;
            16'b1001100011000010: note = 0;
            16'b1001100011010001: note = D1_note;
            16'b1001100101011111: note = 0;
            16'b1001100101101110: note = D1_note;
            16'b1001100111111100: note = 0;
            16'b1001101000001011: note = D1_note;
            16'b1001101010011001: note = 0;
            16'b1001101010101000: note = F1_note;
            16'b1001101100110110: note = 0;
            16'b1001101101000101: note = F1_note;
            16'b1001101111010011: note = 0;
            16'b1001101111100010: note = F1_note;
            16'b1001110001110000: note = 0;
            16'b1001110001111111: note = F1_note;
            16'b1001111000101000: note = 0;
            16'b1001111001010111: note = D1_note;
            16'b1001111011100101: note = 0;
            16'b1001111011110100: note = D1_note;
            16'b1001111110000010: note = 0;
            16'b1001111110010001: note = D1_note;
            16'b1010000000011111: note = 0;
            16'b1010000000101110: note = D1_note;
            16'b1010000010111100: note = 0;
            16'b1010000011001011: note = D1_note;
            16'b1010000101011001: note = 0;
            16'b1010000101101000: note = D1_note;
            16'b1010000111110110: note = 0;
            16'b1010001000000101: note = D1_note;
            16'b1010001010010011: note = 0;
            16'b1010001010100010: note = D1_note;
            16'b1010001100110000: note = 0;
            16'b1010001100111111: note = D1_note;
            16'b1010001111001101: note = 0;
            16'b1010001111011100: note = D1_note;
            16'b1010010001101010: note = 0;
            16'b1010010001111001: note = F1_note;
            16'b1010010100000111: note = 0;
            16'b1010010100010110: note = F1_note;
            16'b1010010110100100: note = 0;
            16'b1010010110110011: note = F1_note;
            16'b1010011001000001: note = 0;
            16'b1010011001010000: note = F1_note;
            16'b1010011111111001: note = 0;
            16'b1010100000101000: note = Dh1_note;
            16'b1010100001101111: note = 0;
            16'b1010100001110111: note = D1_note;
            16'b1010100010111110: note = 0;
            16'b1010100011000110: note = C1_note;
            16'b1010101001101111: note = 0;
            16'b1010101010011110: note = Ah_note;
            16'b1010110101100010: note = 0;
            16'b1010110110110000: note = Ah_note;
            16'b1010111000111110: note = 0;
            16'b1010111001001101: note = F1_note;
            16'b1010111011011011: note = 0;
            16'b1010111011101010: note = F1_note;
            16'b1010111101111000: note = 0;
            16'b1010111110000111: note = F1_note;
            16'b1011000000010101: note = 0;
            16'b1011000000100100: note = F1_note;
            16'b1011000111001101: note = 0;
            16'b1011000111111100: note = Dh1_note;
            16'b1011001001000011: note = 0;
            16'b1011001001001011: note = D1_note;
            16'b1011001010010010: note = 0;
            16'b1011001010011010: note = C1_note;
            16'b1011010001000011: note = 0;
            16'b1011010001110010: note = Ah_note;
            16'b1011010100000000: note = 0;
            16'b1011010100001111: note = C1_note;
            16'b1011100011101110: note = 0;
            16'b1011101111010001: note = D1_note;
            16'b1011110001011111: note = 0;
            16'b1011110001101110: note = D1_note;
            16'b1011110011111100: note = 0;
            16'b1011110100001011: note = D1_note;
            16'b1011110110011001: note = 0;
            16'b1011110110101000: note = D1_note;
            16'b1011111000110110: note = 0;
            16'b1011111001000101: note = D1_note;
            16'b1011111011010011: note = 0;
            16'b1011111011100010: note = D1_note;
            16'b1011111101110000: note = 0;
            16'b1011111101111111: note = D1_note;
            16'b1100000000001101: note = 0;
            16'b1100000000011100: note = D1_note;
            16'b1100000010101010: note = 0;
            16'b1100000010111001: note = D1_note;
            16'b1100000101000111: note = 0;
            16'b1100000101010110: note = D1_note;
            16'b1100000111100100: note = 0;
            16'b1100000111110011: note = F1_note;
            16'b1100001010000001: note = 0;
            16'b1100001010010000: note = F1_note;
            16'b1100001100011110: note = 0;
            16'b1100001100101101: note = F1_note;
            16'b1100001110111011: note = 0;
            16'b1100001111001010: note = F1_note;
            16'b1100010101110011: note = 0;
            16'b1100010110100010: note = D1_note;
            16'b1100011000110000: note = 0;
            16'b1100011000111111: note = D1_note;
            16'b1100011011001101: note = 0;
            16'b1100011011011100: note = D1_note;
            16'b1100011101101010: note = 0;
            16'b1100011101111001: note = D1_note;
            16'b1100100000000111: note = 0;
            16'b1100100000010110: note = D1_note;
            16'b1100100010100100: note = 0;
            16'b1100100010110011: note = D1_note;
            16'b1100100101000001: note = 0;
            16'b1100100101010000: note = D1_note;
            16'b1100100111011110: note = 0;
            16'b1100100111101101: note = D1_note;
            16'b1100101001111011: note = 0;
            16'b1100101010001010: note = D1_note;
            16'b1100101100011000: note = 0;
            16'b1100101100100111: note = D1_note;
            16'b1100101110110101: note = 0;
            16'b1100101111000100: note = F1_note;
            16'b1100110001010010: note = 0;
            16'b1100110001100001: note = F1_note;
            16'b1100110011101111: note = 0;
            16'b1100110011111110: note = F1_note;
            16'b1100110110001100: note = 0;
            16'b1100110110011011: note = F1_note;
            16'b1100111101000100: note = 0;
            16'b1100111101110011: note = Dh1_note;
            16'b1100111110111010: note = 0;
            16'b1100111111000010: note = D1_note;
            16'b1101000000001001: note = 0;
            16'b1101000000010001: note = C1_note;
            16'b1101000110111010: note = 0;
            16'b1101000111101001: note = Ah_note;
            16'b1101010010101101: note = 0;
            16'b1101010011111011: note = Ah_note;
            16'b1101010110001001: note = 0;
            16'b1101010110011000: note = F1_note;
            16'b1101011000100110: note = 0;
            16'b1101011000110101: note = F1_note;
            16'b1101011011000011: note = 0;
            16'b1101011011010010: note = F1_note;
            16'b1101011101100000: note = 0;
            16'b1101011101101111: note = F1_note;
            16'b1101100100011000: note = 0;
            16'b1101100101000111: note = Dh1_note;
            16'b1101100110001110: note = 0;
            16'b1101100110010110: note = D1_note;
            16'b1101100111011101: note = 0;
            16'b1101100111100101: note = C1_note;
            16'b1101101110001110: note = 0;
            16'b1101101110111101: note = Ah_note;
            16'b1101110001001011: note = 0;
            16'b1101110001011010: note = C1_note;
            16'b1110000000111001: note = 0;
            16'b1110101001111011: note = Ah_note;
            16'b1110101100001001: note = 0;
            16'b1110101100011000: note = Ah_note;
            16'b1110101110100110: note = 0;
            16'b1110101110110101: note = Ah_note;
            16'b1110110001000011: note = 0;
            16'b1110110001010010: note = Ah_note;
            16'b1110110011100000: note = 0;
            16'b1110110011101111: note = Ah_note;
            16'b1110110101111101: note = 0;
            16'b1110110110001100: note = Ah_note;
            16'b1110111000011010: note = 0;
            16'b1110111000101001: note = Ah_note;
            16'b1110111010110111: note = 0;
            16'b1110111011000110: note = Ah_note;
            16'b1110111101010100: note = 0;
            16'b1110111101100011: note = Ah_note;
            16'b1110111111110001: note = 0;
            16'b1111000000000000: note = Ah_note;
            16'b1111000010001110: note = 0;
            16'b1111000010011101: note = A_note;
            16'b1111000100101011: note = 0;
            16'b1111000100111010: note = A_note;
            16'b1111000111001000: note = 0;
            16'b1111000111010111: note = A_note;
            16'b1111001001100101: note = 0;
            16'b1111001001110100: note = A_note;
            16'b1111001100000010: note = 0;
            16'b1111001100010001: note = A_note;
            16'b1111010000101100: note = 0;
            16'b1111010001001011: note = Ah_note;
            16'b1111010011011001: note = 0;
            16'b1111010011101000: note = A_note;
            16'b1111010101110110: note = 0;
            16'b1111010110000101: note = G_note;
            16'b1111100111110001: note = 0;
            16'b1111111101011001: note = Ah_note;
            16'b1111111111100111: note = 0;
            16'b1111111111110110: note = Ah_note;
            17'b10000000010000100: note = 0;
            17'b10000000010010011: note = Ah_note;
            17'b10000000100100001: note = 0;
            17'b10000000100110000: note = Ah_note;
            17'b10000000110111110: note = 0;
            17'b10000000111001101: note = Ah_note;
            17'b10000001001011011: note = 0;
            17'b10000001001101010: note = Ah_note;
            17'b10000001011111000: note = 0;
            17'b10000001100000111: note = Ah_note;
            17'b10000001110010101: note = 0;
            17'b10000001110100100: note = Ah_note;
            17'b10000010000110010: note = 0;
            17'b10000010001000001: note = A_note;
            17'b10000010011001111: note = 0;
            17'b10000010011011110: note = A_note;
            17'b10000010101101100: note = 0;
            17'b10000010101111011: note = A_note;
            17'b10000011000001001: note = 0;
            17'b10000011000011000: note = A_note;
            17'b10000011010100110: note = 0;
            17'b10000011010110101: note = A_note;
            17'b10000011111010000: note = 0;
            17'b10000011111101111: note = Ah_note;
            17'b10000100001111101: note = 0;
            17'b10000100010001100: note = A_note;
            17'b10000100100011010: note = 0;
            17'b10000100100101001: note = G_note;
            17'b10000110110010101: note = 0;
            17'b10001001011111101: note = Ah_note;
            17'b10001001110001011: note = 0;
            17'b10001001110011010: note = Ah_note;
            17'b10001010000101000: note = 0;
            17'b10001010000110111: note = Ah_note;
            17'b10001010011000101: note = 0;
            17'b10001010011010100: note = Ah_note;
            17'b10001010101100010: note = 0;
            17'b10001010101110001: note = Ah_note;
            17'b10001010111111111: note = 0;
            17'b10001011000001110: note = Ah_note;
            17'b10001011010011100: note = 0;
            17'b10001011010101011: note = Ah_note;
            17'b10001011100111001: note = 0;
            17'b10001011101001000: note = Ah_note;
            17'b10001011111010110: note = 0;
            17'b10001011111100101: note = A_note;
            17'b10001100001110011: note = 0;
            17'b10001100010000010: note = A_note;
            17'b10001100100010000: note = 0;
            17'b10001100100011111: note = A_note;
            17'b10001100110101101: note = 0;
            17'b10001100110111100: note = A_note;
            17'b10001101001001010: note = 0;
            17'b10001101001011001: note = A_note;
            17'b10001101101110100: note = 0;
            17'b10001101110010011: note = Ah_note;
            17'b10001110000100001: note = 0;
            17'b10001110000110000: note = A_note;
            17'b10001110010111110: note = 0;
            17'b10001110011001101: note = G_note;
            17'b10010000100111001: note = 0;
            17'b10010011010100001: note = Ah_note;
            17'b10010011100101111: note = 0;
            17'b10010011100111110: note = Ah_note;
            17'b10010011111001100: note = 0;
            17'b10010011111011011: note = Ah_note;
            17'b10010100001101001: note = 0;
            17'b10010100001111000: note = Ah_note;
            17'b10010100100000110: note = 0;
            17'b10010100100010101: note = Ah_note;
            17'b10010100110100011: note = 0;
            17'b10010100110110010: note = Ah_note;
            17'b10010101001000000: note = 0;
            17'b10010101001001111: note = Ah_note;
            17'b10010101011011101: note = 0;
            17'b10010101011101100: note = Ah_note;
            17'b10010101101111010: note = 0;
            17'b10010101110001001: note = A_note;
            17'b10010110000010111: note = 0;
            17'b10010110000100110: note = A_note;
            17'b10010110010110100: note = 0;
            17'b10010110011000011: note = A_note;
            17'b10010110101010001: note = 0;
            17'b10010110101100000: note = A_note;
            17'b10010110111101110: note = 0;
            17'b10010110111111101: note = A_note;
            17'b10010111100011000: note = 0;
            17'b10010111100110111: note = Ah_note;
            17'b10010111111000101: note = 0;
            17'b10010111111010100: note = A_note;
            17'b10011000001100010: note = 0;
            17'b10011000001110001: note = G_note;
            17'b10011010011011101: note = 0;
   
        endcase  
    end  
    //лесникК�?Ш
    else if (sw_state == 4'b0101) begin
        case (counter_sec) 
            2'b11: note = A_note;
            8'b10001101: note = 0;
            8'b10011100: note = A_note;
            9'b100101001: note = 0;
            9'b100111000: note = C1_note;
            9'b111000101: note = 0;
            9'b111010100: note = C1_note;
            10'b1001100001: note = 0;
            10'b1001110000: note = D1_note;
            10'b1011111101: note = 0;
            10'b1100001100: note = D1_note;
            10'b1110011001: note = 0;
            10'b1110101000: note = E1_note;
            11'b10000110101: note = 0;
            11'b10001000100: note = E1_note;
            11'b10011010001: note = 0;
            11'b10011100000: note = A_note;
            11'b10101101101: note = 0;
            11'b10101111100: note = A_note;
            11'b11000001001: note = 0;
            11'b11000011000: note = C1_note;
            11'b11010100101: note = 0;
            11'b11010110100: note = C1_note;
            11'b11101000001: note = 0;
            11'b11101010000: note = D1_note;
            11'b11111011101: note = 0;
            11'b11111101100: note = D1_note;
            12'b100001111001: note = 0;
            12'b100010001000: note = E1_note;
            12'b100100010101: note = 0;
            12'b100100100100: note = E1_note;
            12'b100110110001: note = 0;
            12'b100111000000: note = A_note;
            12'b101001001101: note = 0;
            12'b101001011100: note = A_note;
            12'b101011101001: note = 0;
            12'b101011111000: note = C1_note;
            12'b101110000101: note = 0;
            12'b101110010100: note = C1_note;
            12'b110000100001: note = 0;
            12'b110000110000: note = G1_note;
            12'b110010111101: note = 0;
            12'b110011001100: note = G1_note;
            12'b110101011001: note = 0;
            12'b110101101000: note = F1_note;
            12'b110111110101: note = 0;
            12'b111000000100: note = F1_note;
            12'b111010010001: note = 0;
            12'b111010100000: note = A_note;
            12'b111100101101: note = 0;
            12'b111100111100: note = A_note;
            12'b111111001001: note = 0;
            12'b111111011000: note = C1_note;
            13'b1000001100101: note = 0;
            13'b1000001110100: note = C1_note;
            13'b1000100000001: note = 0;
            13'b1000100010000: note = G1_note;
            13'b1000110011101: note = 0;
            13'b1000110101100: note = G1_note;
            13'b1001000111001: note = 0;
            13'b1001001001000: note = F1_note;
            13'b1001011010101: note = 0;
            13'b1001011100100: note = F1_note;
            13'b1001101110001: note = 0;
            13'b1001110000000: note = G1_note;
            13'b1010000001101: note = 0;
            13'b1010000011100: note = G1_note;
            13'b1010010101001: note = 0;
            13'b1010010111000: note = F1_note;
            13'b1010101000101: note = 0;
            13'b1010101010100: note = F1_note;
            13'b1010111100001: note = 0;
            13'b1010111110000: note = E1_note;
            13'b1011001111101: note = 0;
            13'b1011010001100: note = E1_note;
            13'b1011100011001: note = 0;
            13'b1011100101000: note = D1_note;
            13'b1011110110101: note = 0;
            13'b1011111000100: note = D1_note;
            13'b1100001010001: note = 0;
            13'b1100001100000: note = G1_note;
            13'b1100011101101: note = 0;
            13'b1100011111100: note = G1_note;
            13'b1100110001001: note = 0;
            13'b1100110011000: note = F1_note;
            13'b1101000100101: note = 0;
            13'b1101000110100: note = F1_note;
            13'b1101011000001: note = 0;
            13'b1101011010000: note = E1_note;
            13'b1101101011101: note = 0;
            13'b1101101101100: note = E1_note;
            13'b1101111111001: note = 0;
            13'b1110000001000: note = D1_note;
            13'b1110010010101: note = 0;
            13'b1110010100100: note = D1_note;
            13'b1110100110001: note = 0;
            13'b1110101000000: note = G_note;
            13'b1110111001101: note = 0;
            13'b1110111011100: note = G_note;
            13'b1111001101001: note = 0;
            13'b1111001111000: note = B_note;
            13'b1111100000101: note = 0;
            13'b1111100010100: note = B_note;
            13'b1111110100001: note = 0;
            13'b1111110110000: note = C1_note;
            14'b10000000111101: note = 0;
            14'b10000001001100: note = C1_note;
            14'b10000011011001: note = 0;
            14'b10000011101000: note = D1_note;
            14'b10000101110101: note = 0;
            14'b10000110000100: note = D1_note;
            14'b10001000010001: note = 0;
            14'b10001000100000: note = G_note;
            14'b10001010101101: note = 0;
            14'b10001010111100: note = G_note;
            14'b10001101001001: note = 0;
            14'b10001101011000: note = B_note;
            14'b10001111100101: note = 0;
            14'b10001111110100: note = B_note;
            14'b10010010000001: note = 0;
            14'b10010010010000: note = C1_note;
            14'b10010100011101: note = 0;
            14'b10010100101100: note = C1_note;
            14'b10010110111001: note = 0;
            14'b10010111001000: note = D1_note;
            14'b10011001010101: note = 0;
            14'b10011001100100: note = D1_note;
            14'b10011011110001: note = 0;
            14'b10011100000000: note = A_note;
            14'b10011110001101: note = 0;
            14'b10011110011100: note = A_note;
            14'b10100000101001: note = 0;
            14'b10100000111000: note = C1_note;
            14'b10100011000101: note = 0;
            14'b10100011010100: note = C1_note;
            14'b10100101100001: note = 0;
            14'b10100101110000: note = D1_note;
            14'b10100111111101: note = 0;
            14'b10101000001100: note = D1_note;
            14'b10101010011001: note = 0;
            14'b10101010101000: note = E1_note;
            14'b10101100110101: note = 0;
            14'b10101101000100: note = E1_note;
            14'b10101111010001: note = 0;
            14'b10101111100000: note = A_note;
            14'b10110001101101: note = 0;
            14'b10110001111100: note = A_note;
            14'b10110100001001: note = 0;
            14'b10110100011000: note = C1_note;
            14'b10110110100101: note = 0;
            14'b10110110110100: note = C1_note;
            14'b10111001000001: note = 0;
            14'b10111001010000: note = D1_note;
            14'b10111011011101: note = 0;
            14'b10111011101100: note = D1_note;
            14'b10111101111001: note = 0;
            14'b10111110001000: note = E1_note;
            14'b11000000010101: note = 0;
            14'b11000000100100: note = E1_note;
            14'b11000010110001: note = 0;
            14'b11000011000000: note = A_note;
            14'b11000101001101: note = 0;
            14'b11000101011100: note = A_note;
            14'b11000111101001: note = 0;
            14'b11000111111000: note = C1_note;
            14'b11001010000101: note = 0;
            14'b11001010010100: note = C1_note;
            14'b11001100100001: note = 0;
            14'b11001100110000: note = G1_note;
            14'b11001110111101: note = 0;
            14'b11001111001100: note = G1_note;
            14'b11010001011001: note = 0;
            14'b11010001101000: note = F1_note;
            14'b11010011110101: note = 0;
            14'b11010100000100: note = F1_note;
            14'b11010110010001: note = 0;
            14'b11010110100000: note = A_note;
            14'b11011000101101: note = 0;
            14'b11011000111100: note = A_note;
            14'b11011011001001: note = 0;
            14'b11011011011000: note = C1_note;
            14'b11011101100101: note = 0;
            14'b11011101110100: note = C1_note;
            14'b11100000000001: note = 0;
            14'b11100000010000: note = G1_note;
            14'b11100010011101: note = 0;
            14'b11100010101100: note = G1_note;
            14'b11100100111001: note = 0;
            14'b11100101001000: note = F1_note;
            14'b11100111010101: note = 0;
            14'b11100111100100: note = F1_note;
            14'b11101001110001: note = 0;
            14'b11101010000000: note = G1_note;
            14'b11101100001101: note = 0;
            14'b11101100011100: note = G1_note;
            14'b11101110101001: note = 0;
            14'b11101110111000: note = F1_note;
            14'b11110001000101: note = 0;
            14'b11110001010100: note = F1_note;
            14'b11110011100001: note = 0;
            14'b11110011110000: note = E1_note;
            14'b11110101111101: note = 0;
            14'b11110110001100: note = E1_note;
            14'b11111000011001: note = 0;
            14'b11111000101000: note = D1_note;
            14'b11111010110101: note = 0;
            14'b11111011000100: note = D1_note;
            14'b11111101010001: note = 0;
            14'b11111101100000: note = G1_note;
            14'b11111111101101: note = 0;
            14'b11111111111100: note = G1_note;
            15'b100000010001001: note = 0;
            15'b100000010011000: note = F1_note;
            15'b100000100100101: note = 0;
            15'b100000100110100: note = F1_note;
            15'b100000111000001: note = 0;
            15'b100000111010000: note = E1_note;
            15'b100001001011101: note = 0;
            15'b100001001101100: note = E1_note;
            15'b100001011111001: note = 0;
            15'b100001100001000: note = D1_note;
            15'b100001110010101: note = 0;
            15'b100001110100100: note = D1_note;
            15'b100010000110001: note = 0;
            15'b100010001000000: note = G_note;
            15'b100010011001101: note = 0;
            15'b100010011011100: note = G_note;
            15'b100010101101001: note = 0;
            15'b100010101111000: note = B_note;
            15'b100011000000101: note = 0;
            15'b100011000010100: note = B_note;
            15'b100011010100001: note = 0;
            15'b100011010110000: note = C1_note;
            15'b100011100111101: note = 0;
            15'b100011101001100: note = C1_note;
            15'b100011111011001: note = 0;
            15'b100011111101000: note = D1_note;
            15'b100100001110101: note = 0;
            15'b100100010000100: note = D1_note;
            15'b100100100010001: note = 0;
            15'b100100100100000: note = G_note;
            15'b100101000111001: note = 0;
            15'b100101001011000: note = B_note;
            15'b100101101110001: note = 0;
            15'b100101110010000: note = C1_note;
            15'b100110010101001: note = 0;
            15'b100110011001000: note = D1_note;
            15'b100110111100001: note = 0;
            15'b100111000000000: note = A_note;
            15'b100111100011001: note = 0;
            15'b100111100111000: note = C1_note;
            15'b101000001010001: note = 0;
            15'b101000001110000: note = D1_note;
            15'b101000110001001: note = 0;
            15'b101000110101000: note = E1_note;
            15'b101001000110101: note = 0;
            15'b101001001000100: note = A_note;
            15'b101001011010001: note = 0;
            15'b101001101111100: note = A_note;
            15'b101010000001001: note = 0;
            15'b101010000011000: note = C1_note;
            15'b101010100110001: note = 0;
            15'b101010101010000: note = D1_note;
            15'b101011001101001: note = 0;
            15'b101011010001000: note = E1_note;
            15'b101011110100001: note = 0;
            15'b101011111000000: note = A_note;
            15'b101100011011001: note = 0;
            15'b101100011111000: note = C1_note;
            15'b101101000010001: note = 0;
            15'b101101000110000: note = G1_note;
            15'b101101101001001: note = 0;
            15'b101101101101000: note = F1_note;
            15'b101101111110101: note = 0;
            15'b101110000000100: note = A_note;
            15'b101110010010001: note = 0;
            15'b101110100111100: note = A_note;
            15'b101110111001001: note = 0;
            15'b101110111011000: note = C1_note;
            15'b101111011110001: note = 0;
            15'b101111100010000: note = G1_note;
            15'b110000000101001: note = 0;
            15'b110000001001000: note = F1_note;
            15'b110000101100001: note = 0;
            15'b110000110000000: note = G1_note;
            15'b110001010011001: note = 0;
            15'b110001010111000: note = F1_note;
            15'b110001111010001: note = 0;
            15'b110001111110000: note = E1_note;
            15'b110010100001001: note = 0;
            15'b110010100101000: note = D1_note;
            15'b110010110110101: note = 0;
            15'b110010111000100: note = G1_note;
            15'b110011001010001: note = 0;
            15'b110011011111100: note = G1_note;
            15'b110011110001001: note = 0;
            15'b110011110011000: note = F1_note;
            15'b110100010110001: note = 0;
            15'b110100011010000: note = E1_note;
            15'b110100111101001: note = 0;
            15'b110101000001000: note = D1_note;
            15'b110101100100001: note = 0;
            15'b110101101000000: note = G_note;
            15'b110110001011001: note = 0;
            15'b110110001111000: note = B_note;
            15'b110110110010001: note = 0;
            15'b110110110110000: note = C1_note;
            15'b110111011001001: note = 0;
            15'b110111011101000: note = D1_note;
            15'b110111101110101: note = 0;
            15'b110111110000100: note = G_note;
            15'b111000000010001: note = 0;
            15'b111000010111100: note = G_note;
            15'b111000101001001: note = 0;
            15'b111000101011000: note = B_note;
            15'b111001001110001: note = 0;
            15'b111001010010000: note = C1_note;
            15'b111001110101001: note = 0;
            15'b111001111001000: note = D1_note;
            15'b111010011100001: note = 0;
            15'b111010100000000: note = A_note;
            15'b111011000011001: note = 0;
            15'b111011000111000: note = C1_note;
            15'b111011101010001: note = 0;
            15'b111011101110000: note = D1_note;
            15'b111100010001001: note = 0;
            15'b111100010101000: note = E1_note;
            15'b111100100110101: note = 0;
            15'b111100101000100: note = A_note;
            15'b111100111010001: note = 0;
            15'b111101001111100: note = A_note;
            15'b111101100001001: note = 0;
            15'b111101100011000: note = C1_note;
            15'b111110000110001: note = 0;
            15'b111110001010000: note = D1_note;
            15'b111110101101001: note = 0;
            15'b111110110001000: note = E1_note;
            15'b111111010100001: note = 0;
            15'b111111011000000: note = A_note;
            15'b111111111011001: note = 0;
            15'b111111111111000: note = C1_note;
            16'b1000000100010001: note = 0;
            16'b1000000100110000: note = G1_note;
            16'b1000001001001001: note = 0;
            16'b1000001001101000: note = F1_note;
            16'b1000001011110101: note = 0;
            16'b1000001100000100: note = A_note;
            16'b1000001110010001: note = 0;
            16'b1000010000111100: note = A_note;
            16'b1000010011001001: note = 0;
            16'b1000010011011000: note = C1_note;
            16'b1000010111110001: note = 0;
            16'b1000011000010000: note = G1_note;
            16'b1000011100101001: note = 0;
            16'b1000011101001000: note = F1_note;
            16'b1000100001100001: note = 0;
            16'b1000100010000000: note = G1_note;
            16'b1000100110011001: note = 0;
            16'b1000100110111000: note = F1_note;
            16'b1000101011010001: note = 0;
            16'b1000101011110000: note = E1_note;
            16'b1000110000001001: note = 0;
            16'b1000110000101000: note = D1_note;
            16'b1000110010110101: note = 0;
            16'b1000110011000100: note = G1_note;
            16'b1000110101010001: note = 0;
            16'b1000110111111100: note = G1_note;
            16'b1000111010001001: note = 0;
            16'b1000111010011000: note = F1_note;
            16'b1000111110110001: note = 0;
            16'b1000111111010000: note = E1_note;
            16'b1001000011101001: note = 0;
            16'b1001000100001000: note = D1_note;
            16'b1001001000100001: note = 0;
            16'b1001001001000000: note = G_note;
            16'b1001001101011001: note = 0;
            16'b1001001101111000: note = B_note;
            16'b1001010010010001: note = 0;
            16'b1001010010110000: note = C1_note;
            16'b1001010111001001: note = 0;
            16'b1001010111101000: note = D1_note;
            16'b1001011001110101: note = 0;
            16'b1001011010000100: note = G_note;
            16'b1001011100010001: note = 0;
            16'b1001011110111100: note = G_note;
            16'b1001100001001001: note = 0;
            16'b1001100001011000: note = B_note;
            16'b1001100101110001: note = 0;
            16'b1001100110010000: note = C1_note;
            16'b1001101010101001: note = 0;
            16'b1001101011001000: note = D1_note;
            16'b1001101111100001: note = 0;
            16'b1111100011000110: note = A_note;
            16'b1111100101010011: note = 0;
            16'b1111100101100010: note = A_note;
            16'b1111100111101111: note = 0;
            16'b1111100111111110: note = C1_note;
            16'b1111101010001011: note = 0;
            16'b1111101010011010: note = C1_note;
            16'b1111101100100111: note = 0;
            16'b1111101100110110: note = D1_note;
            16'b1111101111000011: note = 0;
            16'b1111101111010010: note = D1_note;
            16'b1111110001011111: note = 0;
            16'b1111110001101110: note = E1_note;
            16'b1111110011111011: note = 0;
            16'b1111110100001010: note = E1_note;
            16'b1111110110010111: note = 0;
            16'b1111110110100110: note = A_note;
            16'b1111111000110011: note = 0;
            16'b1111111001000010: note = A_note;
            16'b1111111011001111: note = 0;
            16'b1111111011011110: note = C1_note;
            16'b1111111101101011: note = 0;
            16'b1111111101111010: note = C1_note;
            17'b10000000000000111: note = 0;
            17'b10000000000010110: note = D1_note;
            17'b10000000010100011: note = 0;
            17'b10000000010110010: note = D1_note;
            17'b10000000100111111: note = 0;
            17'b10000000101001110: note = E1_note;
            17'b10000000111011011: note = 0;
            17'b10000000111101010: note = E1_note;
            17'b10000001001110111: note = 0;
            17'b10000001010000110: note = A_note;
            17'b10000001100010011: note = 0;
            17'b10000001100100010: note = A_note;
            17'b10000001110101111: note = 0;
            17'b10000001110111110: note = C1_note;
            17'b10000010001001011: note = 0;
            17'b10000010001011010: note = C1_note;
            17'b10000010011100111: note = 0;
            17'b10000010011110110: note = G1_note;
            17'b10000010110000011: note = 0;
            17'b10000010110010010: note = G1_note;
            17'b10000011000011111: note = 0;
            17'b10000011000101110: note = F1_note;
            17'b10000011010111011: note = 0;
            17'b10000011011001010: note = F1_note;
            17'b10000011101010111: note = 0;
            17'b10000011101100110: note = A_note;
            17'b10000011111110011: note = 0;
            17'b10000100000000010: note = A_note;
            17'b10000100010001111: note = 0;
            17'b10000100010011110: note = C1_note;
            17'b10000100100101011: note = 0;
            17'b10000100100111010: note = C1_note;
            17'b10000100111000111: note = 0;
            17'b10000100111010110: note = G1_note;
            17'b10000101001100011: note = 0;
            17'b10000101001110010: note = G1_note;
            17'b10000101011111111: note = 0;
            17'b10000101100001110: note = F1_note;
            17'b10000101110011011: note = 0;
            17'b10000101110101010: note = F1_note;
            17'b10000110000110111: note = 0;
            17'b10000110001000110: note = G1_note;
            17'b10000110011010011: note = 0;
            17'b10000110011100010: note = G1_note;
            17'b10000110101101111: note = 0;
            17'b10000110101111110: note = F1_note;
            17'b10000111000001011: note = 0;
            17'b10000111000011010: note = F1_note;
            17'b10000111010100111: note = 0;
            17'b10000111010110110: note = E1_note;
            17'b10000111101000011: note = 0;
            17'b10000111101010010: note = E1_note;
            17'b10000111111011111: note = 0;
            17'b10000111111101110: note = D1_note;
            17'b10001000001111011: note = 0;
            17'b10001000010001010: note = D1_note;
            17'b10001000100010111: note = 0;
            17'b10001000100100110: note = G1_note;
            17'b10001000110110011: note = 0;
            17'b10001000111000010: note = G1_note;
            17'b10001001001001111: note = 0;
            17'b10001001001011110: note = F1_note;
            17'b10001001011101011: note = 0;
            17'b10001001011111010: note = F1_note;
            17'b10001001110000111: note = 0;
            17'b10001001110010110: note = E1_note;
            17'b10001010000100011: note = 0;
            17'b10001010000110010: note = E1_note;
            17'b10001010010111111: note = 0;
            17'b10001010011001110: note = D1_note;
            17'b10001010101011011: note = 0;
            17'b10001010101101010: note = D1_note;
            17'b10001010111110111: note = 0;
            17'b10001011000000110: note = G_note;
            17'b10001011010010011: note = 0;
            17'b10001011010100010: note = G_note;
            17'b10001011100101111: note = 0;
            17'b10001011100111110: note = B_note;
            17'b10001011111001011: note = 0;
            17'b10001011111011010: note = B_note;
            17'b10001100001100111: note = 0;
            17'b10001100001110110: note = C1_note;
            17'b10001100100000011: note = 0;
            17'b10001100100010010: note = C1_note;
            17'b10001100110011111: note = 0;
            17'b10001100110101110: note = D1_note;
            17'b10001101000111011: note = 0;
            17'b10001101001001010: note = D1_note;
            17'b10001101011010111: note = 0;
            17'b10001101011100110: note = G_note;
            17'b10001101111111111: note = 0;
            17'b10001110000011110: note = B_note;
            17'b10001110100110111: note = 0;
            17'b10001110101010110: note = C1_note;
            17'b10001111001101111: note = 0;
            17'b10001111010001110: note = D1_note;
            17'b10001111110100111: note = 0;
            17'b10001111111000110: note = A_note;
            17'b10010000011011111: note = 0;
            17'b10010000011111110: note = C1_note;
            17'b10010001000010111: note = 0;
            17'b10010001000110110: note = D1_note;
            17'b10010001101001111: note = 0;
            17'b10010001101101110: note = E1_note;
            17'b10010001111111011: note = 0;
            17'b10010010000001010: note = A_note;
            17'b10010010010010111: note = 0;
            17'b10010010101000010: note = A_note;
            17'b10010010111001111: note = 0;
            17'b10010010111011110: note = C1_note;
            17'b10010011011110111: note = 0;
            17'b10010011100010110: note = D1_note;
            17'b10010100000101111: note = 0;
            17'b10010100001001110: note = E1_note;
            17'b10010100101100111: note = 0;
            17'b10010100110000110: note = A_note;
            17'b10010101010011111: note = 0;
            17'b10010101010111110: note = C1_note;
            17'b10010101111010111: note = 0;
            17'b10010101111110110: note = G1_note;
            17'b10010110100001111: note = 0;
            17'b10010110100101110: note = F1_note;
            17'b10010110110111011: note = 0;
            17'b10010110111001010: note = A_note;
            17'b10010111001010111: note = 0;
            17'b10010111100000010: note = A_note;
            17'b10010111110001111: note = 0;
            17'b10010111110011110: note = C1_note;
            17'b10011000010110111: note = 0;
            17'b10011000011010110: note = G1_note;
            17'b10011000111101111: note = 0;
            17'b10011001000001110: note = F1_note;
            17'b10011001100100111: note = 0;
            17'b10011001101000110: note = G1_note;
            17'b10011010001011111: note = 0;
            17'b10011010001111110: note = F1_note;
            17'b10011010110010111: note = 0;
            17'b10011010110110110: note = E1_note;
            17'b10011011011001111: note = 0;
            17'b10011011011101110: note = D1_note;
            17'b10011011101111011: note = 0;
            17'b10011011110001010: note = G1_note;
            17'b10011100000010111: note = 0;
            17'b10011100011000010: note = G1_note;
            17'b10011100101001111: note = 0;
            17'b10011100101011110: note = F1_note;
            17'b10011101001110111: note = 0;
            17'b10011101010010110: note = E1_note;
            17'b10011101110101111: note = 0;
            17'b10011101111001110: note = D1_note;
            17'b10011110011100111: note = 0;
            17'b10011110100000110: note = G_note;
            17'b10011111000011111: note = 0;
            17'b10011111000111110: note = B_note;
            17'b10011111101010111: note = 0;
            17'b10011111101110110: note = C1_note;
            17'b10100000010001111: note = 0;
            17'b10100000010101110: note = D1_note;
            17'b10100000100111011: note = 0;
            17'b10100000101001010: note = G_note;
            17'b10100000111010111: note = 0;
            17'b10100001010000010: note = G_note;
            17'b10100001100001111: note = 0;
            17'b10100001100011110: note = B_note;
            17'b10100010000110111: note = 0;
            17'b10100010001010110: note = C1_note;
            17'b10100010101101111: note = 0;
            17'b10100010110001110: note = D1_note;
            17'b10100011010100111: note = 0;
            17'b11000011001000000: note = A_note;
            17'b11000011011001101: note = 0;
            17'b11000011011011100: note = A_note;
            17'b11000011101101001: note = 0;
            17'b11000011101111000: note = C1_note;
            17'b11000100000000101: note = 0;
            17'b11000100000010100: note = C1_note;
            17'b11000100010100001: note = 0;
            17'b11000100010110000: note = D1_note;
            17'b11000100100111101: note = 0;
            17'b11000100101001100: note = D1_note;
            17'b11000100111011001: note = 0;
            17'b11000100111101000: note = E1_note;
            17'b11000101001110101: note = 0;
            17'b11000101010000100: note = E1_note;
            17'b11000101100010001: note = 0;
            17'b11000101100100000: note = A_note;
            17'b11000101110101101: note = 0;
            17'b11000101110111100: note = A_note;
            17'b11000110001001001: note = 0;
            17'b11000110001011000: note = C1_note;
            17'b11000110011100101: note = 0;
            17'b11000110011110100: note = C1_note;
            17'b11000110110000001: note = 0;
            17'b11000110110010000: note = D1_note;
            17'b11000111000011101: note = 0;
            17'b11000111000101100: note = D1_note;
            17'b11000111010111001: note = 0;
            17'b11000111011001000: note = E1_note;
            17'b11000111101010101: note = 0;
            17'b11000111101100100: note = E1_note;
            17'b11000111111110001: note = 0;
            17'b11001000000000000: note = A_note;
            17'b11001000010001101: note = 0;
            17'b11001000010011100: note = A_note;
            17'b11001000100101001: note = 0;
            17'b11001000100111000: note = C1_note;
            17'b11001000111000101: note = 0;
            17'b11001000111010100: note = C1_note;
            17'b11001001001100001: note = 0;
            17'b11001001001110000: note = G1_note;
            17'b11001001011111101: note = 0;
            17'b11001001100001100: note = G1_note;
            17'b11001001110011001: note = 0;
            17'b11001001110101000: note = F1_note;
            17'b11001010000110101: note = 0;
            17'b11001010001000100: note = F1_note;
            17'b11001010011010001: note = 0;
            17'b11001010011100000: note = A_note;
            17'b11001010101101101: note = 0;
            17'b11001010101111100: note = A_note;
            17'b11001011000001001: note = 0;
            17'b11001011000011000: note = C1_note;
            17'b11001011010100101: note = 0;
            17'b11001011010110100: note = C1_note;
            17'b11001011101000001: note = 0;
            17'b11001011101010000: note = G1_note;
            17'b11001011111011101: note = 0;
            17'b11001011111101100: note = G1_note;
            17'b11001100001111001: note = 0;
            17'b11001100010001000: note = F1_note;
            17'b11001100100010101: note = 0;
            17'b11001100100100100: note = F1_note;
            17'b11001100110110001: note = 0;
            17'b11001100111000000: note = G1_note;
            17'b11001101001001101: note = 0;
            17'b11001101001011100: note = G1_note;
            17'b11001101011101001: note = 0;
            17'b11001101011111000: note = F1_note;
            17'b11001101110000101: note = 0;
            17'b11001101110010100: note = F1_note;
            17'b11001110000100001: note = 0;
            17'b11001110000110000: note = E1_note;
            17'b11001110010111101: note = 0;
            17'b11001110011001100: note = E1_note;
            17'b11001110101011001: note = 0;
            17'b11001110101101000: note = D1_note;
            17'b11001110111110101: note = 0;
            17'b11001111000000100: note = D1_note;
            17'b11001111010010001: note = 0;
            17'b11001111010100000: note = G1_note;
            17'b11001111100101101: note = 0;
            17'b11001111100111100: note = G1_note;
            17'b11001111111001001: note = 0;
            17'b11001111111011000: note = F1_note;
            17'b11010000001100101: note = 0;
            17'b11010000001110100: note = F1_note;
            17'b11010000100000001: note = 0;
            17'b11010000100010000: note = E1_note;
            17'b11010000110011101: note = 0;
            17'b11010000110101100: note = E1_note;
            17'b11010001000111001: note = 0;
            17'b11010001001001000: note = D1_note;
            17'b11010001011010101: note = 0;
            17'b11010001011100100: note = D1_note;
            17'b11010001101110001: note = 0;
            17'b11010001110000000: note = G_note;
            17'b11010010000001101: note = 0;
            17'b11010010000011100: note = G_note;
            17'b11010010010101001: note = 0;
            17'b11010010010111000: note = B_note;
            17'b11010010101000101: note = 0;
            17'b11010010101010100: note = B_note;
            17'b11010010111100001: note = 0;
            17'b11010010111110000: note = C1_note;
            17'b11010011001111101: note = 0;
            17'b11010011010001100: note = C1_note;
            17'b11010011100011001: note = 0;
            17'b11010011100101000: note = D1_note;
            17'b11010011110110101: note = 0;
            17'b11010011111000100: note = D1_note;
            17'b11010100001010001: note = 0;
            17'b11010100001100000: note = G_note;
            17'b11010100101111001: note = 0;
            17'b11010100110011000: note = B_note;
            17'b11010101010110001: note = 0;
            17'b11010101011010000: note = C1_note;
            17'b11010101111101001: note = 0;
            17'b11010110000001000: note = D1_note;
            17'b11010110100100001: note = 0;
            17'b11010110101000000: note = A_note;
            17'b11010111001011001: note = 0;
            17'b11010111001111000: note = C1_note;
            17'b11010111110010001: note = 0;
            17'b11010111110110000: note = D1_note;
            17'b11011000011001001: note = 0;
            17'b11011000011101000: note = E1_note;
            17'b11011000101110101: note = 0;
            17'b11011000110000100: note = A_note;
            17'b11011001000010001: note = 0;
            17'b11011001010111100: note = A_note;
            17'b11011001101001001: note = 0;
            17'b11011001101011000: note = C1_note;
            17'b11011010001110001: note = 0;
            17'b11011010010010000: note = D1_note;
            17'b11011010110101001: note = 0;
            17'b11011010111001000: note = E1_note;
            17'b11011011011100001: note = 0;
            17'b11011011100000000: note = A_note;
            17'b11011100000011001: note = 0;
            17'b11011100000111000: note = C1_note;
            17'b11011100101010001: note = 0;
            17'b11011100101110000: note = G1_note;
            17'b11011101010001001: note = 0;
            17'b11011101010101000: note = F1_note;
            17'b11011101100110101: note = 0;
            17'b11011101101000100: note = A_note;
            17'b11011101111010001: note = 0;
            17'b11011110001111100: note = A_note;
            17'b11011110100001001: note = 0;
            17'b11011110100011000: note = C1_note;
            17'b11011111000110001: note = 0;
            17'b11011111001010000: note = G1_note;
            17'b11011111101101001: note = 0;
            17'b11011111110001000: note = F1_note;
            17'b11100000010100001: note = 0;
            17'b11100000011000000: note = G1_note;
            17'b11100000111011001: note = 0;
            17'b11100000111111000: note = F1_note;
            17'b11100001100010001: note = 0;
            17'b11100001100110000: note = E1_note;
            17'b11100010001001001: note = 0;
            17'b11100010001101000: note = D1_note;
            17'b11100010011110101: note = 0;
            17'b11100010100000100: note = G1_note;
            17'b11100010110010001: note = 0;
            17'b11100011000111100: note = G1_note;
            17'b11100011011001001: note = 0;
            17'b11100011011011000: note = F1_note;
            17'b11100011111110001: note = 0;
            17'b11100100000010000: note = E1_note;
            17'b11100100100101001: note = 0;
            17'b11100100101001000: note = D1_note;
            17'b11100101001100001: note = 0;
            17'b11100101010000000: note = G_note;
            17'b11100101110011001: note = 0;
            17'b11100101110111000: note = B_note;
            17'b11100110011010001: note = 0;
            17'b11100110011110000: note = C1_note;
            17'b11100111000001001: note = 0;
            17'b11100111000101000: note = D1_note;
            17'b11100111010110101: note = 0;
            17'b11100111011000100: note = G_note;
            17'b11100111101010001: note = 0;
            17'b11100111111111100: note = G_note;
            17'b11101000010001001: note = 0;
            17'b11101000010011000: note = B_note;
            17'b11101000110110001: note = 0;
            17'b11101000111010000: note = C1_note;
            17'b11101001011101001: note = 0;
            17'b11101001100001000: note = D1_note;
            17'b11101010000100001: note = 0;
            17'b11111101101010000: note = B_note;
            17'b11111110001101001: note = 0;
            17'b11111110010001000: note = D1_note;
            17'b11111110110100001: note = 0;
            17'b11111110111000000: note = E1_note;
            17'b11111111011011001: note = 0;
            17'b11111111011111000: note = Fh1_note;
            17'b11111111110000101: note = 0;
            17'b11111111110010100: note = B_note;
            18'b100000000000100001: note = 0;
            18'b100000000011001100: note = B_note;
            18'b100000000101011001: note = 0;
            18'b100000000101101000: note = D1_note;
            18'b100000001010000001: note = 0;
            18'b100000001010100000: note = E1_note;
            18'b100000001110111001: note = 0;
            18'b100000001111011000: note = Fh1_note;
            18'b100000010011110001: note = 0;
            18'b100000010100010000: note = B_note;
            18'b100000011000101001: note = 0;
            18'b100000011001001000: note = D1_note;
            18'b100000011101100001: note = 0;
            18'b100000011110000000: note = A1_note;
            18'b100000100010011001: note = 0;
            18'b100000100010111000: note = G1_note;
            18'b100000100101000101: note = 0;
            18'b100000100101010100: note = B_note;
            18'b100000100111100001: note = 0;
            18'b100000101010001100: note = B_note;
            18'b100000101100011001: note = 0;
            18'b100000101100101000: note = D1_note;
            18'b100000110001000001: note = 0;
            18'b100000110001100000: note = A1_note;
            18'b100000110101111001: note = 0;
            18'b100000110110011000: note = G1_note;
            18'b100000111010110001: note = 0;
            18'b100000111011010000: note = A1_note;
            18'b100000111111101001: note = 0;
            18'b100001000000001000: note = G1_note;
            18'b100001000100100001: note = 0;
            18'b100001000101000000: note = Fh1_note;
            18'b100001001001011001: note = 0;
            18'b100001001001111000: note = E1_note;
            18'b100001001100000101: note = 0;
            18'b100001001100010100: note = A1_note;
            18'b100001001110100001: note = 0;
            18'b100001010001001100: note = A1_note;
            18'b100001010011011001: note = 0;
            18'b100001010011101000: note = G1_note;
            18'b100001011000000001: note = 0;
            18'b100001011000100000: note = Fh1_note;
            18'b100001011100111001: note = 0;
            18'b100001011101011000: note = E1_note;
            18'b100001100001110001: note = 0;
            18'b100001100010010000: note = A_note;
            18'b100001100110101001: note = 0;
            18'b100001100111001000: note = Ch1_note;
            18'b100001101011100001: note = 0;
            18'b100001101100000000: note = D1_note;
            18'b100001110000011001: note = 0;
            18'b100001110000111000: note = E1_note;
            18'b100001110011000101: note = 0;
            18'b100001110011010100: note = A_note;
            18'b100001110101100001: note = 0;
            18'b100001111000001100: note = A_note;
            18'b100001111010011001: note = 0;
            18'b100001111010101000: note = Ch1_note;
            18'b100001111111000001: note = 0;
            18'b100001111111100000: note = D1_note;
            18'b100010000011111001: note = 0;
            18'b100010000100011000: note = E1_note;
            18'b100010001000110001: note = 0;
            18'b100010001001010000: note = B_note;
            18'b100010001101101001: note = 0;
            18'b100010001110001000: note = D1_note;
            18'b100010010010100001: note = 0;
            18'b100010010011000000: note = E1_note;
            18'b100010010111011001: note = 0;
            18'b100010010111111000: note = Fh1_note;
            18'b100010011010000101: note = 0;
            18'b100010011010010100: note = B_note;
            18'b100010011100100001: note = 0;
            18'b100010011111001100: note = B_note;
            18'b100010100001011001: note = 0;
            18'b100010100001101000: note = D1_note;
            18'b100010100110000001: note = 0;
            18'b100010100110100000: note = E1_note;
            18'b100010101010111001: note = 0;
            18'b100010101011011000: note = Fh1_note;
            18'b100010101111110001: note = 0;
            18'b100010110000010000: note = B_note;
            18'b100010110100101001: note = 0;
            18'b100010110101001000: note = D1_note;
            18'b100010111001100001: note = 0;
            18'b100010111010000000: note = A1_note;
            18'b100010111110011001: note = 0;
            18'b100010111110111000: note = G1_note;
            18'b100011000001000101: note = 0;
            18'b100011000001010100: note = B_note;
            18'b100011000011100001: note = 0;
            18'b100011000110001100: note = B_note;
            18'b100011001000011001: note = 0;
            18'b100011001000101000: note = D1_note;
            18'b100011001101000001: note = 0;
            18'b100011001101100000: note = A1_note;
            18'b100011010001111001: note = 0;
            18'b100011010010011000: note = G1_note;
            18'b100011010110110001: note = 0;
            18'b100011010111010000: note = A1_note;
            18'b100011011011101001: note = 0;
            18'b100011011100001000: note = G1_note;
            18'b100011100000100001: note = 0;
            18'b100011100001000000: note = Fh1_note;
            18'b100011100101011001: note = 0;
            18'b100011100101111000: note = E1_note;
            18'b100011101000000101: note = 0;
            18'b100011101000010100: note = A1_note;
            18'b100011101010100001: note = 0;
            18'b100011101101001100: note = A1_note;
            18'b100011101111011001: note = 0;
            18'b100011101111101000: note = G1_note;
            18'b100011110100000001: note = 0;
            18'b100011110100100000: note = Fh1_note;
            18'b100011111000111001: note = 0;
            18'b100011111001011000: note = E1_note;
            18'b100011111101110001: note = 0;
            18'b100011111110010000: note = A_note;
            18'b100100000010101001: note = 0;
            18'b100100000011001000: note = Ch1_note;
            18'b100100000111100001: note = 0;
            18'b100100001000000000: note = D1_note;
            18'b100100001100011001: note = 0;
            18'b100100001100111000: note = E1_note;
            18'b100100001111000101: note = 0;
            18'b100100001111010100: note = A_note;
            18'b100100010001100001: note = 0;
            18'b100100010100001100: note = A_note;
            18'b100100010110011001: note = 0;
            18'b100100010110101000: note = Ch1_note;
            18'b100100011011000001: note = 0;
            18'b100100011011100000: note = D1_note;
            18'b100100011111111001: note = 0;
            18'b100100100000011000: note = E1_note;
            18'b100100100100110001: note = 0;
            18'b100100110100111000: note = A_note;
            18'b100101000110011101: note = 0;
        endcase  
    end 
    //toxic
    else if (sw_state == 4'b0101) begin
        case (counter_sec) 
            2'b11: note = Ah2_note;
            8'b10010110: note = 0;
            8'b10100111: note = Ah2_note;
            9'b100111101: note = 0;
            9'b101001110: note = Ah2_note;
            9'b111100100: note = 0;
            9'b111110101: note = Ah2_note;
            10'b1010001011: note = 0;
            10'b1010011100: note = B2_note;
            10'b1111001000: note = 0;
            10'b1111101001: note = Gh2_note;
            11'b10100010101: note = 0;
            11'b10100110110: note = Dh3_note;
            11'b11001100010: note = 0;
            11'b11010000011: note = Dh3_note;
            11'b11110101111: note = 0;
            11'b11111010000: note = Ch3_note;
            12'b100011111100: note = 0;
            12'b100100011101: note = B2_note;
            12'b101001001001: note = 0;
            12'b101001101010: note = Ah2_note;
            12'b101110010110: note = 0;
            12'b101110110111: note = Ah2_note;
            12'b110011100011: note = 0;
            12'b110100000100: note = B2_note;
            12'b111000110000: note = 0;
            12'b111001010001: note = Gh2_note;
            12'b111101111101: note = 0;
            12'b111110011110: note = Ah2_note;
            13'b1000011001010: note = 0;
            13'b1000011101011: note = B2_note;
            13'b1001000010111: note = 0;
            13'b1001000111000: note = Ah2_note;
            13'b1001101100100: note = 0;
            13'b1001110000101: note = Gh2_note;
            13'b1010010110001: note = 0;
            13'b1010011010010: note = G2_note;
            13'b1010111111110: note = 0;
            13'b1011000011111: note = G2_note;
            13'b1011101001011: note = 0;
            13'b1011101101100: note = Gh2_note;
            13'b1100010011000: note = 0;
            13'b1100010111001: note = Gh2_note;
            13'b1100111100101: note = 0;
            13'b1101000000110: note = Dh3_note;
            13'b1101100110010: note = 0;
            13'b1101101010011: note = Dh3_note;
            13'b1101111101001: note = 0;
            13'b1101111111010: note = Dh3_note;
            13'b1110010010000: note = 0;
            13'b1110010100001: note = Ch3_note;
            13'b1110111001101: note = 0;
            13'b1110111101110: note = B2_note;
            13'b1111100011010: note = 0;
            13'b1111100111011: note = Ah2_note;
            14'b10000001100111: note = 0;
            14'b10000010001000: note = Ah2_note;
            14'b10000110110100: note = 0;
            14'b10000111010101: note = B2_note;
            14'b10001100000001: note = 0;
            14'b10001100100010: note = Gh2_note;
            14'b10010001001110: note = 0;
            14'b10010001101111: note = Ah2_note;
            14'b10010110011011: note = 0;
            14'b10010110111100: note = B2_note;
            14'b10011011101000: note = 0;
            14'b10011100001001: note = Ah2_note;
            14'b10100000110101: note = 0;
            14'b10100001010110: note = B2_note;
            14'b10100110000010: note = 0;
            14'b10100110100011: note = Ah2_note;
            14'b10101011001111: note = 0;
            14'b10101011110000: note = B2_note;
            14'b10110000011100: note = 0;
            14'b10110000111101: note = Gh2_note;
            14'b10110101101001: note = 0;
        endcase  
    end  
end

endmodule